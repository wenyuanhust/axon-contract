{
  "deployment": {
    "lock": {
      "code_hash": "0x9bd7e06f3ecf4be0f2fcd2188b23f1b9fcc88e5d4b65a8637b17723bbda3cce8",
      "hash_type": "type",
      "args": "0x61a0d1fa2b4a4536a778659d5d87b88e82188b17"
    },
    "cells": [
      {
        "name": "stake",
        "location": {
          "file": "build/release/stake"
        },
        "enable_type_id": true
      },
      {
        "name": "stake-smt",
        "location": {
          "file": "build/release/stake-smt"
        },
        "enable_type_id": true
      }
    ],
    "dep_groups": [],
    "multisig_config": {
      "sighash_addresses": [],
      "require_first_n": 0,
      "threshold": 0
    }
  },
  "last_recipe": null,
  "new_recipe": {
    "cell_recipes": [
      {
        "name": "stake",
        "tx_hash": "0x45a9fd2d766fb0afe0f1003362cfba03aa0a66d4ec5e036c0cdbebe4d9dabcac",
        "index": 0,
        "occupied_capacity": 16298200000000,
        "data_hash": "0xcc8a15b5b0ed1f413a417e5b633bcc2992ef4963c02d86661c8528af10b6074d",
        "type_id": "0x4eb776810a6050036422b4c8e96deb2f75e4a5cb89f598f7d31d282b9e761929"
      },
      {
        "name": "stake-smt",
        "tx_hash": "0x45a9fd2d766fb0afe0f1003362cfba03aa0a66d4ec5e036c0cdbebe4d9dabcac",
        "index": 1,
        "occupied_capacity": 26771000000000,
        "data_hash": "0xb84cc4290ebff4aa996da56cfb3ae1102745f94b136b1c1137c535532a9bfe6f",
        "type_id": "0x2a250a7bd74c42c3c9a56934c93ee9e8b488553325dca476631fd7c96d3728c9"
      }
    ],
    "dep_group_recipes": []
  },
  "used_input_txs": {
    "0x45a9fd2d766fb0afe0f1003362cfba03aa0a66d4ec5e036c0cdbebe4d9dabcac": {
      "version": "0x0",
      "cell_deps": [
        {
          "out_point": {
            "tx_hash": "0xf8de3bb47d055cdf460d93a2a6e1b05f7432f9777c8c474abf4eec1d4aee5d37",
            "index": "0x0"
          },
          "dep_type": "dep_group"
        }
      ],
      "header_deps": [],
      "inputs": [
        {
          "since": "0x0",
          "previous_output": {
            "tx_hash": "0xbe3777fa551ec2de85ece9cca9918eefc953db190d52426d74c5f1cc73b2868c",
            "index": "0x1"
          }
        },
        {
          "since": "0x0",
          "previous_output": {
            "tx_hash": "0xe6a4b80a06bbfbdb23456e6845b8ee87aa9644ad185c25295c919dbe6dbd8da0",
            "index": "0x1"
          }
        }
      ],
      "outputs": [
        {
          "capacity": "0xed2b86be600",
          "lock": {
            "code_hash": "0x9bd7e06f3ecf4be0f2fcd2188b23f1b9fcc88e5d4b65a8637b17723bbda3cce8",
            "hash_type": "type",
            "args": "0x61a0d1fa2b4a4536a778659d5d87b88e82188b17"
          },
          "type": {
            "code_hash": "0x00000000000000000000000000000000000000000000000000545950455f4944",
            "hash_type": "type",
            "args": "0xb7fe83392736c6d1633f35194d1a0e7e87fcc908a84394074031b5b95e06c026"
          }
        },
        {
          "capacity": "0x18591bf1fe00",
          "lock": {
            "code_hash": "0x9bd7e06f3ecf4be0f2fcd2188b23f1b9fcc88e5d4b65a8637b17723bbda3cce8",
            "hash_type": "type",
            "args": "0x61a0d1fa2b4a4536a778659d5d87b88e82188b17"
          },
          "type": {
            "code_hash": "0x00000000000000000000000000000000000000000000000000545950455f4944",
            "hash_type": "type",
            "args": "0xf89735de346f9655e16d60c3d91963fe67f8b845f511e5fcdea60d462c94a33e"
          }
        },
        {
          "capacity": "0x12d9e4a31c3fd",
          "lock": {
            "code_hash": "0x9bd7e06f3ecf4be0f2fcd2188b23f1b9fcc88e5d4b65a8637b17723bbda3cce8",
            "hash_type": "type",
            "args": "0x61a0d1fa2b4a4536a778659d5d87b88e82188b17"
          },
          "type": null
        }
      ],
      "outputs_data": [
        "0x7f454c460201010000000000000000000200f30001000000d426010000000000400000000000000028770200000000000100000040003800050040001400120006000000040000004000000000000000400001000000000040000100000000001801000000000000180100000000000008000000000000000100000004000000000000000000000000000100000000000000010000000000d416000000000000d41600000000000000100000000000000100000005000000d416000000000000d426010000000000d4260100000000001c850000000000001c8500000000000000100000000000000100000006000000f09b000000000000f0bb010000000000f0bb01000000000028010000000000002821080000000000001000000000000051e574640600000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c740100000000005e74010000000000707401000000000088740100000000009e7401000000000020950100000000001e95010000000000229501000000000026950100000000002a95010000000000c874010000000000000000000000000001000000000000003686010000000000617474656d707420746f206164642077697468206f766572666c6f7700000000617474656d707420746f2073756274726163742077697468206f766572666c6f7700000000000000c87401000000000001000000000000000100000000000000088c01000000000008c9bcf367e6096a3ba7ca8485ae67bb2bf894fe72f36e3cf1361d5f3af54fa5d182e6ad7f520e511f6c3e2b8c68059b6bbd41fbabd9831f79217e1319cde05bc874010000000000000000000000000001000000000000000c800100000000000000000000000000617474656d707420746f207368696674206c6566742077697468206f766572666c6f7700000000000000000000000000617474656d707420746f206d756c7469706c792077697468206f766572666c6f77000000000000000000000000000000617474656d707420746f2073756274726163742077697468206f766572666c6f77000000000000000000000000000000617474656d707420746f2073686966742072696768742077697468206f766572666c6f77000000000000000000000000617474656d707420746f206164642077697468206f766572666c6f776c6561662073697a65206d75737420626520616c69676e20746f203136206279746573007c0301000000000023000000000000007265717569726573206d6f7265206d656d6f727920737061636520746f20696e697469616c697a65204275646479416c6c6f630000000000b00301000000000033000000000000006f7574206f66206d656d6f72790000000000000000000000617474656d707420746f20646976696465206279207a65726f00000000000000617474656d707420746f206164642077697468206f766572666c6f77427974655265616465724279746533325265616465724279746573526561646572000000617474656d707420746f2073756274726163742077697468206f766572666c6f775363726970745265616465725769746e65737341726773526561646572556e6b6e6f776e000000c874010000000000080000000000000008000000000000007a88010000000000456e636f64696e674f766572666c6f7776616c69646174654c656e6774684e6f74456e6f75676800c874010000000000080000000000000008000000000000007a880100000000004974656d4d697373696e67496e6465784f75744f66426f756e6429426f72726f774572726f72426f72726f774d75744572726f7200000000787701000000000018000000000000000800000000000000b880010000000000748201000000000028830100000000002020202052656164446174612c0a2c20280a282c30783030303130323033303430353036303730383039313031313132313331343135313631373138313932303231323232333234323532363237323832393330333133323333333433353336333733383339343034313432343334343435343634373438343935303531353235333534353535363537353835393630363136323633363436353636363736383639373037313732373337343735373637373738373938303831383238333834383538363837383838393930393139323933393439353936393739383939000078770100000000000800000000000000080000000000000060830100000000006a8301000000000020840100000000002829000000000000787701000000000008000000000000000800000000000000208601000000000054727946726f6d536c6963654572726f72636b622d64656661756c742d68617368616c726561647920626f72726f77656400000000000000c874010000000000000000000000000001000000000000000c80010000000000616c7265616479206d757461626c7920626f72726f776564c87401000000000000000000000000000100000000000000fa7f01000000000063616c6c656420604f7074696f6e3a3a756e77726170282960206f6e206120604e6f6e65602076616c75650000000000c87401000000000001000000000000000100000000000000088c010000000000617474656d707420746f206164642077697468206f766572666c6f77726561645f6174206069662073697a65203c20726561645f6c656e60726561645f6174206069662064732e63616368655f73697a65203e2064732e6d61785f63616368655f73697a6560726561645f617420606966206375722e6f6666736574203c2064732e73746172745f706f696e74207c7c202e2e2e60726561645f61742060696620726561645f706f696e74202b20726561645f6c656e203e2064732e63616368655f73697a656076616c69646174653a2073697a65203e206375722e736f757263652e746f74616c5f73697a65756e7061636b5f6e756d6265726765745f6974656d5f636f756e74636f6e766572745f746f5f753634636f6e766572745f746f5f7538636f6e7665727420746f205665633c75383e00000096910100000000001800000000000000080000000000000062900100000000004669656c64436f756e744f75744f66426f756e64556e6b6e6f776e4974656d4f6666736574486561646572546f74616c53697a65436f6d6d6f6e0000000000000000000000000000617474656d707420746f206164642077697468206f766572666c6f770000000063616c6c65642060526573756c743a3a756e77726170282960206f6e20616e2060457272602076616c75650000000000c874010000000000000000000000000001000000000000003686010000000000c874010000000000100000000000000008000000000000003674010000000000617373657274696f6e206661696c65643a20636865636b706f696e745f646174612e69735f6e6f6e652829617373657274696f6e206661696c65643a207374616b655f61745f646174612e69735f6e6f6e6528290000000006000000000000000900000000000000060000000000000006000000000000000b000000000000000a000000000000000a000000000000000400000000000000080000000000000004000000000000002c0901000000000023090100000000001d0901000000000017090100000000000c090100000000000209010000000000f8080100000000009005010000000000e0040100000000008c050100000000001000000000000000017a5200017801011b0c02002c00000018000000061c0000181b000000440ed00d74810188028903920493059406950796089709980a990b9a0c9b0d1000000048000000ee3600000a000000000e0000100000005c000000e436000008000000000000001000000070000000d836000008000000000000001c00000084000000cc3600004e00000000420e304a810188028903920493050018000000a4000000fa3600003000000000420e20468101880289030014000000c00000000e3700000e00000000420e104281010014000000d8000000043700000e00000000420e104281010018000000f0000000fa3600005800000000420e404481018802000000180000000c010000363700005800000000420e4044810188020000001800000028010000723700005800000000420e4044810188020000001800000044010000ae3700005800000000420e4044810188020000001400000060010000ea3700005200000000420e40428101001800000078010000243800005800000000420e4044810188020000001400000094010000603800005200000000420e404281010018000000ac0100009a3800005800000000420e40448101880200000018000000c8010000d63800004e00000000420e3044810188020000001c000000e4010000083900009a00000000420e20488101880289039204000000200000000402000082390000dc00000000440e304c8101880289039204930594060000002c000000280200003a3a0000ee1a000000420ef0035a810188028903920493059406950796089709980a990b9a0c9b0d2c00000058020000f85400001404000000420e80015a810188028903920493059406950796089709980a990b9a0c9b0d1000000088020000dc5800003c000000000e0000100000009c020000045900000a000000000e000010000000b0020000fa5800004c000000000e000010000000c4020000325900004c000000000e000010000000d80200006a590000f4000000000e00002c000000ec0200004a5a0000d403000000420eb00158810188028903920493059406950796089709980a990b9a0c00002c0000001c030000ee5d0000f203000000420ec0015a810188028903920493059406950796089709980a990b9a0c9b0d200000004c030000b0610000d600000000420e504e8101880289039204930594069507001800000070030000626200005200000000420e204681018802890300140000008c030000986200003400000000420e104281010018000000a4030000b46200007400000000420e50468101880289030014000000c00300000c6300003600000000420e104281010020000000d80300002a6300006c00000000420e304c81018802890392049305940600000020000000fc030000726300006200000000420e304c8101880289039204930594060000001000000020040000b063000022000000000e00001800000034040000be6300003a00000000420e2046810188028903002000000050040000dc630000fc00000000420e404e8101880289039204930594069507001000000074040000b464000042000000000e00001400000088040000e26400009200000000420e104281010010000000a00400005c650000020000000000000010000000b40400004a650000360000000000000018000000c80400006c6500007a00000000420e40448101880200000018000000e4040000ca6500008200000000420e4044810188020000002400000000050000306600006001000000440ee0086481018802890392049305940695079608970910000000280500006867000018000000000e0000100000003c0500006c670000040000000000000010000000500500005c670000020000000000000014000000640500004a6700004201000000420e30428101002c0000007c05000074680000e401000000420e705a810188028903920493059406950796089709980a990b9a0c9b0d001c000000ac050000286a00005600000000420e304a810188028903920493050024000000cc0500005e6a00007803000000420e50528101880289039204930594069507960897090014000000f4050000ae6d00000e00000000420e1042810100240000000c060000a46d00007e01000000420e8001508101880289039204930594069507960800001000000034060000fa6e000012000000000000001000000048060000f86e00001200000000000000140000005c060000f66e00000e00000000420e10428101001400000074060000ec6e00000e00000000420e1042810100140000008c060000e26e00000e00000000420e104281010014000000a4060000d86e00007000000000420e90014281012c000000bc060000306f0000bc01000000420e90015a810188028903920493059406950796089709980a990b9a0c9b0d14000000ec060000bc700000b400000000420e10428101001400000004070000587100003800000000420e4042810100100000001c070000787100000a0000000000000014000000300700006e710000b600000000420e104281010014000000480700000c7200003a00000000420e404281010020000000600700002e7200002001000000420ea0014e81018802890392049305940695071c000000840700002a7300009800000000420e4048810188028903920400000014000000a4070000a27300000e00000000420e104281010010000000bc07000098730000160000000000000018000000d00700009a730000a200000000420e40468101880289030014000000ec070000207400007000000000420e90014281011c00000004080000787400005200000000420e304a81018802890392049305001800000024080000aa7400007e00000000420e5046810188028903001c000000400800000c7500006200000000420e2048810188028903920400000010000000600800004e750000300000000000000018000000740800006a7500004e00000000420e1044810188020000001c000000900800009c7500006800000000420e304a810188028903920493050018000000b0080000e47500007e00000000420e50468101880289030018000000cc080000467600005200000000420e20468101880289030018000000e80800007c7600005600000000420e1044810188020000002000000004090000b67600008201000000420e504e8101880289039204930594069507001000000028090000147800002800000000000000100000003c090000287800006200000000420e101800000050090000767800006800000000420e304481018802000000180000006c090000c27800005400000000420e3044810188020000002400000088090000fa7800007c01000000420e80015281018802890392049305940695079608970918000000b00900004e7a00007800000000420e40468101880289030018000000cc090000aa7a00007e00000000420e4046810188028903001c000000e80900000c7b0000a200000000420e5048810188028903920400000018000000080a00008e7b00007a00000000420e20468101880289030020000000240a0000ec7b0000ba00000000420e504c81018802890392049305940600000010000000480a0000827c00001000000000000000100000005c0a00007e7c0000080000000000000010000000700a0000727c0000080000000000000010000000840a0000667c0000080000000000000010000000980a00005a7c0000080000000000000010000000ac0a00004e7c00000a000000000e00001c000000c00a0000447c00007200000000420e5048810188028903920400000024000000e00a0000967c0000ca02000000420ea0015081018802890392049305940695079608000010000000080b0000387f000028000000000e0000240000001c0b00004c7f00006401000000420ea0015081018802890392049305940695079608000024000000440b0000888000008605000000440e800864810188028903920493059406950796089709280000006c0b0000e68500001803000000420eb00256810188028903920493059406950796089709980a990b18000000980b0000d28800009200000000420eb001468101880289032c000000b40b000048890000a003000000420ed0025a810188028903920493059406950796089709980a990b9a0c9b0d24000000e40b0000b88c00008601000000420e90014c8101880289039204930594060000000000000000000002452c00014697000000e78000019308d00573000000130101932334116c2330816c233c916a2338216b2334316b2330416b233c5169233861692334716923308169233c91672338a1672334b167179600001306665e0ce208e6080c1306004013040040814597800000e78040db2338816205659b08458093050163080c09440146814601478147014873000000aa84630285080545638da406114463900418033b01631305004063786507854505445a8597600000e7804012aa8cae8a0c0c1306004097800000e78040e293020bc013850c402338516285659b88458093050163130600400943814601478147014873000000630d6510aa846309851011446397041083340163094463e29210a1a0014429a2054419a25a85814597600000e780a00baa8cae8a0c0c5a8697800000e780c0db114463708b023145b14b814597600000e78060092a892e8a17e5ffff930515c791a003c51c0083c50c0003c62c0083c63c0022054d8d4206e206558e3364a600631a8b02214463788b0e3145b14b814597600000e78020052a892e8a17e5ffff9305d5c231464a8597800000e780c0d485442da03145b14b814597600000e78080022a892e8a17e5ffff930535c031464a8597800000e78020d28144da8923289120232a8121233c8120233031232334212323384123233c7123080c97500000e78060c00d4463870a00668597700000e780a08dda8409a8014463870a00668597700000e780608c2285a68597700000e78080c12a841315840361958330816c0334016c8334816b0339016b8339816a033a016a833a8169033b0169833b8168033c0168833c8167033d0167833d81661301016d828003c55c0083c54c0003c66c0083c67c0022054d8d4206e206558e3364a6001335840093753400b335b0004d8d15c531453149814597600000e78080f32a84ae8917e5ffff930535b13146228597800000e78020c38d4409bf63708b023145b14b814597600000e780a0f02a892e8a17e5ffff930555ae65bd93592400fd190d4563f8a9023145b14b814597600000e78020ee2a892e8a17e5ffff9305d5ab31464a8597800000e780c0bd91440d446dbd639ea908114691446685da85a28697500000e780008a13f63500f199b306b5002338a120233cb1202330d1222334c12223389122130501630c0c97400000e780005a13050163da8597500000e7808088033901638334016423382121233c912009452330a122080c97500000e780e09921cd31453149814597600000e78040e42a84ae8917e5ffff9305f5a13146228597800000e780e0b38d4459aa3145b14b814597600000e780a0e12a892e8a17e5ffff9305559f31464a8597800000e78040b10d449144cdbb6380047605456380a47603360900833689006685da8597400000e780007d13040002639e850e09456382a47403368900833609016685da8597400000e780e07a0544639e850e0d456385a47203360901833689016685da8597400000e780e0782a86ae86080cb285368697400000e780807d8324012115456393a4100335816311c54a8597600000e78040672d45636465016f10e00d93054bff0d456364b5006f10c00403c5dc0083c5cc0003c6ec0083c6fc0022054d8d4206e206558e83c51c0083c60c0003c72c0083873c00a205d58d4207e2075d8fd98d1147b366a600638ce50a03c55c0083c54c0003c66c0003877c0022054d8d42066207598e518d8d4563f6a56a7199c1456317b508080ce6855a8697400000e78000674da8ae893145b14b814597600000e780e0cc2a892e8a17e5ffff9305e586314605a0ae892945a94b814597600000e780e0ca2a892e8a17e5ffff9305458429464a8597800000e780809a814403358163e30205c80335016397600000e780405895b9032c4121033481218339012203398122033a0123833b8123c9bf93050bff0d45e377b57403c51c0183c50c0103c62c0103c73c0122054d8d42066207598e3367a600080ce6855a8697400000e78020550334012103360122281a9146a28597400000e780805a0335812111c5228597600000e780c0507279b6642685814597600000e78080bf2a84ae89ca85268697800000e780a08f23388120233c312123309122130501630c0c97600000e780004003390163033481631305016313070002ca852286814697600000e780000003350163e30405720335016483358163033601632330a122233cb1202338c120880a0c0c97600000e780a02913050163930600025147ca85228697600000e780e0fb03350163e30c056e0335016483358163033601632330a122233cb1202338c120a8120c0c97600000e7808025080c1306004013040040814597700000e78020772338816205659b08a581054562151307150093050163080c01468146814701487300000021c54944567511c5367597600000e780c03f766511c5566597600000e780e03e4a8597600000e78060c6166511c5727597600000e780603de38f0ab0668597600000e780803c01be033a0163130510406367aa0685450544528597600000e78080aaaa892efa0c0c1306004097700000e780807a93040ac0138509402338916285659b88a581131784030507930501631306004081468147014873000000833501633335a000b3b5b4004d8d21c9527529d94e8597600000e780203599b75285814597600000e78000a4aa892efa0c0c528697700000e7802074114463708a024545454c814597600000e780c0a12a8bae8b17d5ffff9305356091a003c5190083c5090003c6290083c6390022054d8d4206e206558e3364a600631a8a02214463788a084545454c814597600000e780809d2a8bae8b17d5ffff9305f55b45465a8597700000e780206d054d2da04545454c814597600000e780e09a2a8bae8b17d5ffff9305555945465a8597700000e780806a014d2328a121232ab121233c8120233041232334612323387123233c8123080c97400000e780e05849445275e30205e64e8597600000e780002699bd03c5590083c5490003c6690083c6790022054d8d4206e206558e3364a6001335840093753400b335b0004d8d15c54545454b814597600000e780e0912a842e8a17d5ffff930555504546228597700000e78080610d4d85bf63708a024545454c814597600000e780008f2a8bae8b17d5ffff9305754d21bf93542400fd140d4563f8a4024545454c814597600000e780808c2a8bae8b17d5ffff9305f54a45465a8597700000e780205c114d0d44e1a0639ea408114691444e85d285a28697400000e780602813f63500f199b306b5002338a120233cb1202330d1222334c12223389122130501630c0c97400000e78060f813050163d28597400000e780e026033b01630334016423386121233c812009452330a122080c97400000e780403829cd4545454b814597600000e780a0822a842e8a17d5ffff930515414546228597700000e78040520d4d75a24545454c814597600000e78000802a8bae8b17d5ffff9305753e45465a8597700000e780a04f0d44114d268ab9b56302041405456302a41403360b0083368b004e85d28597400000e780401b99cd2a86ae86080cb285368697400000e780c01f032d012115456316ad1209456309a41003368b0083360b014e85d28597400000e780c01799cd2a86ae86080cb285368697400000e780401c032d01211545631aad0e0d456300a40e03360b0183368b014e85d28597400000e780401499cd2a86ae86080cb285368697400000e780c018032d01211545631ead0a0335816311c55a8597600000e780800293058aff0d45e377b52093054affe373b52003c5990083c5890003c6a90083c6b90022054d8d4206e206558eb366a60003c5d90083c5c90003c6e90003c7f90022054d8d42066207598e3367a600080cce85528697400000e780c0fe033501222aee49c503340121f2642685814597500000e780e06a2a8a2eeaa285268697700000e780003ba5a00145814509a80545854531a00945894519a00d458d4597500000e780603e0000832d412103348121033a0122033b8122833b0123033c812303358163e30605cc0335016397600000e78040f575b917d5ffff1305c5209305100297500000e780e0bf0000014a0335812119c50335012197600000e78080f263080a3a0d45f265e37cb55a03451a0083450a0003462a0083063a0022054d8d4206e206558e518d854529446318b554167593050002e31fb568d667014b02f603c5970183c5870103c6a70183c6b70122054d8d4206e206558e518d83c5d70103c6c70183c6e70103c7f701a205d18dc2066207d98ed58d82154d8daae303c5170183c5070103c6270183c6370122054d8d4206e206558e518d83c5570103c6470183c6670103c77701a205d18dc2066207d98ed58d82154d8d2aff03c5970083c5870003c6a70083c6b70022054d8d4206e206558e518d83c5d70003c6c70083c6e70003c7f700a205d18dc2066207d98ed58d82154d8d2afb03c5170083c5070003c6270083c6370022054d8d4206e206558e518d83c5570003c6470083c667003ee603c77700a205d18dc2066207d98ed58d82154d8d2af70d45aaff23300120130d1121930d9165080cac1b97600000e78040df034501218945630cb5246303051003459d0183458d010346ad018346bd0122054d8d4206e206558e518d8345dd010346cd018346ed010347fd01a205d18dc2066207d98ed58d82154d8d2334a16403451d0183450d0103462d0183463d0122054d8d4206e206558e518d83455d0103464d0183466d0103477d01a205d18dc2066207d98ed58d82154d8d2330a16403459d0083458d000346ad008346bd0022054d8d4206e206558e518d8345dd000346cd008346ed000347fd00a205d18dc2066207d98ed58d82154d8d233ca16203451d0083450d0003462d0083463d0022054d8d4206e206558e518d83455d0003464d0083466d0003477d00a205d18dc2066207d98ed58d82154d8d2338a16209a82334016423300164233c016223380162130501632c131306000297700000e780604d012519c1b27419aa130501630d46da8597400000e780600d03340163e301042e033581632af2833401642685814597500000e7806036aa8b2e8ca285268697700000e780800623387163233c816323309164130501659305016397600000e780c0b60385ed008385dd0003c6cd0083340165230fa162a205d18d231eb16203c59d0083c58d0003c6ad008386bd0022054d8d4206e206558e518d232ca16203c51d0083c50d0003c62d0083c63d0022054d8d4206e20683c55d00558e518d03c64d00a20583c66d0003c77d00d18d834b8165c2066207d98ed58d82154d8d2338a162327511c5327597500000e78020430305e1638315c16303268163833601632307a11e2316b11e2324c11eb6f3127511c5228597600000e78040b87d556300ab56050b26f671bb294419b232756301051c0305e11e8315c11e0326811e9e76230ba11c231ab11c2328c11cb6e713051162ac033d4697700000e78000f53275233ca16023007163080c930581610d4697500000e780806c033b0121e3010b2e0305712283056122034651222303a11aa205d18d2312b11a0345212283451122034631228306412222054d8d4206e206558e518d2320a11a0345a121834591210346b1218346c12122054d8d4206e2068345e121558e518d0346d121a2058346f12103470122d18d03048121c2066207d98ed58d82154d8d2aef327597500000e780e031130591182c0b3d4697700000e780a0e95ae323048118130501630c030d4697500000e780606103350163e30505240335016483358163033601632330a122233cb1202338c12028130c0c97600000e780c085130501630c03114697500000e780a05d03350163e30005220335016483358163033601632330a122233cb1202338c120130501630c0c97600000e780e081ba7d7a768334016303370164080cee85a68697600000e780c0ed0c0c13060002326597700000e7808021833581632a8491c5268597600000e780009d5a7511c56e8597600000e780209c0dc45a8597500000e78080231304300319a01304b0065265630d05f2528597600000e780c0996ff0cff2080c9146d285726697400000e78040a1833b0121833401222685814597500000e78000072a842e8bde85268697700000e78020d7e38004168344040063070b00228597600000e780e0940335812119c50335012197600000e780c093526511c5528597600000e780e0920545638aa4024944639b042e080c0546814597400000e78060c60345012163090510033581218335012297600000e780a0c52a84e9a4130501650c0397100000e780a0af28130c0397100000e780e0a3130501630c0397100000e78080a83a747a768334016303370164080ca285a68697600000e78000da13050002814597500000e78040faaa8b2e8b0c0c1306000297700000e78040ca0335816311c5268597600000e78060885a7511c5228597600000e780808793050002054685445e8597700000e78000a21375f50f13043004631e95029305000209465e8597700000e78040a01375f50f13044004631095028334016583350166268597600000e78020bb2a841375f50f630c052063070b005e8597600000e7804081033581656300051e0335016597600000e7800080c1aa0305712183056121034651212307a11aa205d18d2316b11a0345212183451121034631218306412122054d8d4206e206558e518d2324a11a033581228305012303348121833401222338a162230cb1621305f11b93050163254697700000e780a0ba13558403230ba11a13550403a30aa11a13558402230aa11a13550402a309a11a135584012309a11a13550401a308a11a135584002308a11aa307811a13d58403230fa11a13d50403a30ea11a13d58402230ea11a13d50402a30da11a13d58401230da11a13d50401a30ca11a13d58400230ca11aa30b911a130501650c0397100000e780a0a7080c0c0397100000e78020810334016503360166833401210337012213050163a285a68697600000e78040bd0335812111c5268597500000e780a06d0335816511c5228597500000e780a06c13050002814597500000e78080dbaa8d2e8b930501631306000297700000e78060aba8030c0397100000e780c08a3e65fe6597600000e78060a12a841375f50f05ed080cac03054697600000e78020400345012105e10334812283340122080cac03094697600000e780603e0345012163020510034411215e6511c53e6597500000e780406463070b006e8597500000e78060631375f40f29c11a6597500000e78080ea6ff06fbb17d5ffff1305c5daf1456ff02fed11456ff08fe863070b005e8597500000e78000600335816511c5268597500000e780005f1a6597500000e78080e6527511c54e8597500000e780805d567511c5367597500000e780a05c766511c5566597500000e780c05b4a8597500000e78040e3166511c5727597500000e780405a63870a00668597500000e780605901446fe0dfcd3145da856ff02fe017d5ffff130525d397c5ffff9386255e09a817d5ffff130505d297c5ffff9386055d9305b002100c97400000e780803c00000335012283358122258da18d4d8d3d44e31a05ee080c2c13054697600000e780e034833b012263880b0c033581212af60335812283350123033681238336012136f22338a164233cb1642330c166aefbaaf7def3080c2c13094697600000e780e030033c0122630b0c08033581212aee0335812283350123033681238336012136ea2338a164233cb1642330c1662334b1202330a120e2ff881397000000e780c0719374f50fa81b97000000e780e0701375f50f51446399a43c130501658c1397000000e780207f080cac1b97000000e780607e03360166033501226313a602833501210335016597700000e780c0c9133a150001a80344012129b50344012149ae014a0335812119c50335012197500000e78000440335816519c50335016597500000e780e04263000a36130581618c1397000000e780807d080c9305816197000000e780806c8335012241456397a54403350121834585002ee583459500aefc8345a500aef88345b500aef48345c500aef08345d5002efc8345e5002ef88345f5002ef4834505002ee183451500aeec83452500aee883453500aee483454500aee0834555002ef0834565002eec833581210346750032e889c597500000e78020391305816197000000e780e05e2ae613050165ac1b97000000e7802073080c9305016597000000e78020628335012241456394a53a03350121834585002ee2834495008345a500aef98345b500aef58345c500aef18345d5002ef98345e5002ef58345f5002ef183450500aefd83451500aeed83452500aee983453500aee583454500aee1834555002eed834565002ee983358121034a750089c597500000e780002f1305016597000000e780c0542afd1305016597000000e780805e2a8d080c13060002ee8597600000e78040d30345012101c503441121d1aa8335812113852500636eb52a130460036311ad1c4a752205aa75c2050a7662066a682208ca68c208620a939284004e7342032e7462048e76b363d500d18d6e6e220ece66c2062e6762070e65b367a800b3641a01126533e5a20033646400b3e575006e763366ce00d98ec58f418d8215558e8217b3e8a50033e8c7000346811085428347810b6315560a62762206c276c206a274e2048273a20362634203c26ee20e667f220f467e420e267a620a0675b36fa600c58ee660a200466d420da665e205066533e7a30033e66e002a653364af003365ca01b3e6f6018a64b3e49000b3e5a501598e418d8216c58d0216c98e4d8e639857043337c800ba876384d800b3b7d8006395071c3275f265638aa50e3275f265c5a817d5ffff1305c59497d5ffff938645999305b002130601652db1639457083275f2656380a5023275f26531a83275f2656383a5043275f26589a01145f2656ff0af9d1275d26533b6a500631d0616127652673335c700b275f266b385b640898d3305c740b3c5b8003345a8004d8d1304700329e56da01275d2653337b500631907141277d26433359700b275f2679d8d898d33059740b58d318d4d8d1304a00311ed32756386a80032753335150121a01275333505011304800335c10335016597500000e780c0950335816197500000e7800095628597500000e78060945e8597500000e780c093a5b41275d265b3b7a500ede73385d840198db305c84012775266b334e600b276f267b386d740858e198e358db18d4d8d1304900345f10335016597500000e780a08f0335816197500000e780e08e628597500000e780408e5e8597500000e780a08d014411b417c5ffff1305e57f97c5ffff93866504f9bc17c5ffff1305c57e97c5ffff9386c5099305b00213060163e9b417c5ffff1305257d97c5ffff938625084dbc17c5ffff1305057c97c5ffff9386050745b417c5ffff1305e5599305b0026ff02f8b17c5ffff1305e500c9ba17c5ffff130545026ff08f8917c5ffff130585016ff0cf8817c5ffff1305c5006ff00f8817c5ffff130505006ff04f8741456ff0ef8297300000e780a0550000172300006700635f173300006700239c797106f422f026ec4ae84ee43284ae892a89328597200000e780205daa8405c163e38900a2892685ca854e8697600000e78040374a8597300000e78040982685a2700274e2644269a26945618280011106ec22e826e42a8497200000e780e058aa8401c926858145228697600000e78080262685e2604264a26405618280411106e497400000e780c0d90000411106e497400000e780e0d80000397106fc22f82a840a85194697500000e780c0a802650dc14265a26502662af42ef032ec2c08228597500000e78020cee27042742161828017c5ffff1305256797c5ffff938625f29305b002300897400000e780a0d10000397106fc22f82a840a851d4697500000e78040a302650dc14265a26502662af42ef032ec2c08228597500000e780a0c8e27042742161828017c5ffff1305a56197c5ffff9386a5ec9305b002300897400000e78020cc0000397106fc22f82a840a85214697500000e780c09d02650dc14265a26502662af42ef032ec2c08228597500000e78020c3e27042742161828017c5ffff1305255c97c5ffff938625e79305b002300897400000e780a0c60000397106fc22f82a840a85354697500000e780409802650dc14265a26502662af42ef032ec2c08228597500000e780a0bde27042742161828017c5ffff1305a55697c5ffff9386a5e19305b002300897400000e78020c10000397106fcaa852800014697500000e780e092226519cd6265c26522662af82ef432f0081097500000e78080b0e2702161828017c5ffff1305855197c5ffff938685dc9305b002101097400000e78000bc0000397106fc22f82a840a85054697500000e780a08d02650dc14265a26502662af42ef032ec2c08228597500000e78000b3e27042742161828017c5ffff1305054c97c5ffff938605d79305b002300897400000e78080b60000397106fcaa852800094697500000e7804088226519cd6265c26522662af82ef432f0081097500000e780609ee2702161828017c5ffff1305e54697c5ffff9386e5d19305b002101097400000e78060b10000397106fc22f82a840a85154697500000e780008302650dc14265a26502662af42ef032ec2c08228597500000e78060a8e27042742161828017c5ffff1305654197c5ffff938665cc9305b002300897400000e780e0ab0000797106f422f02a840a85194697400000e780807d026519c94265a265026608e80ce410e0a27002744561828017c5ffff1305a53c97c5ffff9386a5c79305b0021306f10197400000e78000a70000011106ec22e826e44ae02e892a84130505041306800b814597600000e780e0f117c5ffff930505c613060004228597600000e78060fd13053900a14522868346e5ff0347d5ff8347f5ff83440500a206d98ec207e204c58f0347150083442500dd8e834735000217a214458fc217830445005d8f1c62d98ee214c58ebd8e14e2fd1521062105c5fd0345090068f4e2604264a26402690561828069ce797106f422f026ec4ae84ee452e03284ae842a89687193050008b389a54063f6c9082330090e130a09065295a6854e8697600000e78060380335090493050508033689042330b904133505f81345150032952334a9044a85d28597000000e78000083304344113051008ce94636fa402930900080335090493050508033689042330b904133505f81345150032952334a9044a85a68597000000e7804004130404f893840408e3e789fc0335090e4a9513050506a685228697600000e780e02f0335090e22952330a90ea2700274e2644269a269026a45618280417186f7a2f3a6efcaebcee7d2e356ff5afb5ef762f366ef6aeb6ee72e892a842801130600082401814597600000e78060d90d0941458345e9ff0346d9ff8346f9ff03470900a205d18dc206620703461900d98e03472900d58d0216834639002217598e03074900c216558ed18d6217d98d8ce07d15a104210955fd280213060004a28597600000e780a0e02c603064833204053267b2772a65aae89776000083b46642033884053e972a97a58db98d9774000083b4a44193d605028215d58d338e9500b346fe004a652ae193d78601a216dd8e2a973303d700b345b30013d70501c215b3e8e500469eb345de0093d6f50386055267d274ea67bee4177500000335653db3ebd50026973e97318d398d9775000083b5a53c135605020215518daa95ad8c8a7636f813d68401a214d18c3386e600330996003345a900935605014215b36cd500338abc0033459a009355f5030605f26672772a769774000083b48438b369b500ba96b296328c32f433c59200358d9774000083b464379357050202155d8daa94258fca752eec935787012217d98fae96b382f60033c5a200935605014215b36dd500ee94a58f13d5f703860792761666ea75aefc177700000337873333eba700b296ae963345e800358d177700000337a7329355050202154d8d2a97398e8e67bef0935586012216d18dbe96b383b60033c5a300135605014215518d2a97b98dae6a13d6f5038605d18d56934e933345a300135605020215498eb29433c53401ce69935685012215c98e338569004ee8b30ed50033c6ce00935706014216336df600b3009d0033c6d0006e6f9356f6030606b36fd6007a99fae033032b01b347130193d407028217c58f3e97b34467010e75aaf493d88401a21433e61401b3086500b298b3c7f80093d40701c21733e39700330be3003346cb002e75aaf81357f6030606b364e600aa92ae9233c69201135706020216598e329eb345be004e7913d78501a2154d8fb30559004af03388e5003346c800935206014216b36256003386c201318fee751355f7030607336ea700ae93ae86aeecde9333c5b301935d050202153365b501b30c4501b3cd7c01926793d58d01a21db3e5bd00be933e873efcb38db30033c5ad00935305014215336a750033059a01a98d93d7f5038605dd8db69eae9eb3c76e0093d607028217dd8e3696b18d93d78501a215dd8db387ee01b38eb700b3c6de0093d70601c216b3e3f6003383c300b345b30013d6f5038605b3ecc500e298fe98b3c5120113d605028215d18d2e953346f501935686012216d18e56e4338658013696b18d93d70501c215b3e8f500b382a80033c5d2009355f50306054d8d4e982698b3450a0193d605028215cd8eb690b3c5900093d78501a215cd8fb3050701b38ff500b3c6df0093d40601c21633e89600c290b3c6f00093d7f6038606d58fca9df29db3c6ad0193d406028216d58c338f6401b346cf0113d78601a216558fe676ee96338ae600b3449a0093d50401c214c58d2e9f3347ef009354f7030607d98c8a66b69eaa9eb3c5be0013d705028215d98d33871500398d935685012215c98e467b33856e01b30ed500b3c5be0013d50501c215b3eba500338deb00b346dd0013d5f6038606b3e0a600466c62963e96334576009355050202154d8d2a9fb345ff0093d68501a215d58d266e7296b309b60033c5a900935605014215558d2a9fb345bf0093d6f5038605b3edd5002676b29fa69fb3c51f0193d605028215cd8e3693b345930093d48501a215cd8c8675fe95b3839500b3c6d30093d70601c216d58f3e93b346930093d4f6038606b3e8960062673a9a669ab3460a0193d406028216c58eb692b3c4920193d58401a214c58d4279b3044901b38fb400b3c6df0093d40601c21633ea9600b3045a00a58d93d6f5038605d58db29eae9e33c5ae00935605020215c98eb382660033c5b200935585012215c98d33855e01b30cb500b3c6dc0013d50601c216b3eea600f69233c5b2009355f50306053363b50033063b010696b18f13d5070282175d8d3388a400b345180093d68501a215d58d62962e96318d935605014215b360d50006983345b8009355f50306054d8dba93ee93b3457a0093d605028215cd8eb387a601b3c5b70113d78501a215b3e4e500b385c301338a9500b346da0013d70601c216b3e3e6009e97bd8c93d6f4038604c58ee275ae9fc69fb3c47f0113d704028214458f3a9fb3441f0193d58401a214c58d827bde9fae9f33c7ef00935407014217458f3a9fb345bf0093d4f503860533ec95008665ae9caa9c33c7ec00935407020217458fba973d8d935485012215c98ce669338599012695298f935807014217336b1701b30cfb0033c79c009357f7030607b36df700ca8a4a96b305d60033c7be009357070202175d8fb307ef00bd8e93d48601a216c58e66762e96338dc6003346ed00135706014216b36ee600338efe00b346de0013d7f603860633efe6000676329a629a33471a00935407020217458fba92b3c5820193d48501a215cd8c8a68b3854801338a95003347ea00935707014217336cf700e292b3c7920093d4f7038607b3e097004267ba9f9a9fb3c77f0093d407028217c58f3e98b344680093d68401a214c58e2279ca9fb69fb3c7ff0093d50701c217dd8db3870501bd8e93d4f6038606c58e329536953346d501935406020216458e33085600b346d80093d48601a216c58e3a953695298e935406014216336396001a983346d8009356f6030606b362d600569d6e9d3346ac01935606020216d18eb69733c6b701135786012216598e3387a801b30ac700b3c6da0093d40601c216b3e39600b38df30033c6cd009356f6030606558e5e9a7a9ab3c5450193d605028215cd8eb3889601b3c5e80193d78501a215cd8fc675d295338ab700b346da0093d40601c21633ef9600fa98b3c7f80093d4f7038607c58fa675ae9f869fb3c66f0193d406028216d58cb38ec401b3c61e0093d58601a216d58db3863f01b38fb600b3c49f0093d60401c214c58eb69eb3c5be0093d4f5038605c58da66b5e953307c500b98e93d406028216c58eb69833c6c800935486012216458e66753a953295a98e93d40601c21633ec9600b30c1c0133c6cc009356f6030606336ed600e26833871a013e9733466700935606020216558e3303d601b346f30093d78601a216dd8e866a5697330dd7003346cd00135706014216598e3293b346d30013d7f6038606b3e0e600ca894a9a2e9ab3467a0013d706028216d98e3698b345b80013d78501a215d98dc66433079a00b38ee500b3c6de0093d70601c216dd8e3698b345b80093d7f5038605b3e3f5006279ca9f969fb3c5ef0193d705028215cd8fbe9db3c55d0013d78501a2154d8f226bb305fb01338fe500b347ff0093d50701c217dd8dae9d33c7ed009357f70306075d8fc2673e953a95298e9357060202165d8e32983347e8009357870122175d8f2695b307e5003d8e135506014216b362a60016983345e8001356f5030605518d2ae8469d729d33c5a601135605020215498eb29d33c5cd01935685012215c98e06756a95330dd5003346cd00135706014216b36fe600338ebf013346de009356f6030606d18ede9e869eb3c5d50113d605028215d18db388950133c61800135786012216598e33873e01b30dc700b3c5bd0093d40501c215b3ee9500f698b3c5c80013d6f50386054d8e569f1e9fb3458f0193d405028215cd8c2693b345730013d58501a2154d8db3052f01b383a500b3c4930093d50401c214c58db3846500258d1357f5030605498f6665aa97b697bd8d13d5050282154d8daa98b3c5d80093d68501a215d58d8a66be96b380b60033c5a000935705014215336af500b30b1a0133c5bb009355f50306053363b50026794a9d329d33c5a201935505020215c98db388b40033c5c800135685012215498e467c33058d01330fc500b345bf0093d70501c215cd8fbe98b3c5c80013d6f5038605b3e2c500667dea9dba9db3c5fd0113d605028215d18d2e983346e800135786012216518f33866d01da89b30ce600b3c5bc0093d40501c215c58d2e983347e8009354f7030607b36f9700c27dee934265aa9333c7d301935407020217d98cb38ac40133c7aa00135587012217598d027e33077e00b30ea700b3c49e0013d60401c214d18c33865401318d9356f5030605558da666b690aa90b3c6f00093d706028216dd8eb38a060133c5aa009357850122155d8db3878001aa97bd8e13d70601c21633e8e600c29a33c5aa009356f5030605b363d5006a9f1a9f33c5e501935505020215c98d2e9633456600935685012215c98e06657a95330dd500b345bd0013d70501c21533e3e500330fc300b345df0013d6f5038605d18d4665aa9c969c33c69401935606020216558eb29bb3c65b0013d78601a216558fb3862c013309d7003346c900935406014216336b9600da9b33c6eb001357f6030606598ece9efe9e33c74e01935407020217d98ca69833c7f801935687012217d98e3387be01330cd700b3449c0013d70401c214458fb3041701a58e13d5f6038606c98e2275aa97ae973d8f135507020217598db30f7501b3c5bf0013d78501a215d98df297338ab7003345aa00135705014215b362e500969f33c5bf008e689355f5030605b369b500469d329d33450d019355050202154d8db30e950033c6ce00ca7d135786012216598eb384ad01338dc4003345ad00135705014215498fba9e33c6ce00926c9357f6030606b36bf60066993699334669009357060202165d8eb29ab3c6da0093d78601a216dd8ee667ca97338ed7003346ce00135506014216518daa9a33c6da009356f60306063369d6008a652e9c1e9c33468b01935606020216d18e369f33467f004e68935786012216d18f33060c01338bc700b346db0013d60601c216558eb306e601b58fae7493d5f7038607dd8dd294ae94258f9357070202175d8f330f5701b3c5e50193d78501a215cd8fb385b401338cb70033478701935407014217336a9700529f33c7e701ca679354f703060733639700ea97ce973d8d135705020215598db303d500b3c6790013d78601a216558fb3869701b30cd70033459501935705014215b369f500ce93334577006e779357f50306055d8d72975e97398e9357060202165d8eb29fb3c7fb014e7e93d48701a217c58f7297338de7003346a601135706014216b36ae600d69f33c6f7012a779357f60306065d8e5a974a97b3c5e20093d705028215cd8fbe9eb345d901ee6693d48501a215cd8cb305d700b382b400b3c7570093d60701c217dd8eb69e33c7d401aa679354f7030607d98ce297aa97bd8e13d706028216d98eb69f3345f501135785012215598dc697330cf500b3c6860113d70601c21633e9e6004ae3ca9f3345f501ea761357f5030605b36be500e696b2963345da00135705020215598d330ad501334646018a7e135786012216598ef696b30dd6003345b501935605014215558d2a9a334646019356f6030606336bd600429d269d33c6a901935606020216558e329fb3c6e401ea6493d58601a216d58db3069d00b38cd50033469601935406014216458e329fb3c5e501ae6493d7f5038605b3e9f500a6929a92b3c55a0093d705028215cd8fbe93b34573008e7493d68501a215cd8eb3859200b38ab600b3c7570193d50701c217dd8db3877500bd8e13d7f6038606d98e629e369e3345c501135705020215598db302e501b3c6560013d78601a216d98e269e338cc60133458501135705014215b363e5009e9233c556009356f5030605336fd5007af6ee98de9833451601135605020215518d3303f50033c66b00ee76135786012216598ec696b30bd60033457501935605014215336ed5007293334566002e769356f5030605558d66965a96b18d93d605028215d58db386f5013347db00ca67935487012217d98c3e96338bc400b3c5650113d60501c215b3efc500fe96b58c93d5f4038604b3ecb400d69ece9eb345d90113d605028215d18d2e9a33c64901935486012216d18c33860e01b38ac400b3c5550113d60501c215d18d2e9a33c64401ca741357f6030606598ee294aa94a58d13d705028215d98dae96358d2a679357850122155d8d2697330de500b3c5a50113d70501c215b3eee50076e3b388de0033451501126c9356f50306053369d500e29be69b33c57301935605020215c98eb383460133c57c002a77935785012215c98f3385eb00338aa700b3c6460113d70601c216558fba93b3c677002e6893d7f6038606b3ebf600429b329bb3466e0193d706028216d58fbe9233465600ea75935686012216558eb306bb00330bd600b3c7670113d50701c2175d8daa92334656006a6e9357f6030606b369f600f29afa9a33c65f01935706020216d18f3e9333466f00ee66935486012216d18c3386da002696b18f93d60701c217dd8e3693b3c7640093d4f7038607c58fea95be952d8f935407020217d98ca69233c75700935787012217d98fe295b38ab700b3c4540193d50401c214b3efb400fe92b3c5570093d7f503ee74860533eff5007af6d294ca94258d935505020215c98d2e9333456900ce67135785012215498f3385f400330ca700b3c5850193d70501c21533eaf5005293b34567000e7793d7f5038605cd8f5a975e97b98e93d506028216d58dae98b3c61b018a7413d58601a216558d2697b304e500a58d93d60501c21533e9d500ca9833451501aa659356f5030605558db295ce9533c6be00935606020216558eb293b3c6790013d78601a216d98ec2953388b60033460601135706014216598eb293b3c676002e7793d5f6038606d58d56973e97398e935606020216558eb298b3c6170193d78601a216d58fb306c701b389d70033463601135706014216b36ee60076e3f69833c617014e779357f6030606336bf60062972a9733c6ef00935706020216d18fbe93334575008e6f135685012215518d3306f701330cc500b3c7870113d70701c2175d8fba93334575004a6e9357f5030605b36af500f294ae9433459a009357050202155d8daa92b3c555002a7a13d68501a215d18dd294b38c950033459501135605014215336dc500ea92b3c555006e6693d6f5038605b3ebd50032987a98b345090193d605028215cd8eb3846600b3459f004a7393d78501a215cd8fb30568003389b700b3c6260193d50601c216d58dae94a58f93d6f7038607dd8e4e963696318f9357070202175d8f33085700b3c60601ea6713d58601a216558d3e96b30dc5003347b701135607014217b369c7004e98334505011356f5032e670605336fc5007af662975a973345ed00135605020215518db302950033465b009357860122165d8e5297330be60033456501135705014215336ae500d292334556001356f5030605518de69fd69fb3c5f50113d605028215d18d3387150133c6ea00ea74935786012216d18f33869f00b38fc700b3c5f50193d40501c215b3e895004697b98f93d5f7038607dd8d4a9e5e9eb3c7ce0193d407028217c58fbe93b3c47b0013d68401a214458e7293b30e6600b3c7d70193d40701c217c58fbe933346760092649356f6030606558eee94aa94a58f93d607028217dd8e3383e600334565000e779357850122155d8d2697b30be500b3c6760193d70601c21633eef60072e3729333456500ce669357f50306053369f500da96ae9633c5d900935705020215c98fbe9333c57500ee75935485012215c98c3385b600338ba400b3c7670193d50701c217dd8dae93b3c674008a7a93d7f6038606b3e9f600d69fb29fb346fa0193d706028216dd8e369833460601ae77935486012216458efe97330cf600b3c6860193d40601c216c58e369833460601ce741355f6030606336aa600a69efa9e33c5d801135605020215518daa9233465f002a67935486012216458eba9e330fd6013345e5019357050142155d8daa92334656009357f60306065d8e5e973297b98d93d705028215dd8d2e9833460601ca67935486012216d18c3306f700b38cc400b3c5950113d70501c215b3efe5007e98b3c5040113d7f503ea678605b3eee50076f6da97ca97bd8e93d506028216cd8eb3885600b345190113d78501a2154d8fb3855701330bb700b3c6660193d70601c216b3eaf600d69833471701aa779354f7030607458fe297ce973d8d935405020215458d2a93b3c46900ca7693d58401a214c58dbe96b38bd500334575019356050142153369d5004a9333c56500ea759356f5030605c98efa95d2953345be00935405020215c98ca69333457a008e67135685012215498e3385f500330ca600b3c4840193d50401c214c58db38775003d8eae629354f6030606458e969cba9cb3c5950193d405028215c58db3836500334777004e63935487012217458fb3846c00330d9700b3c5a50113d50501c21533efa500fa9333457700ee6c9355f5030605b369b500669b369b33c56f019355050202154d8daa97bd8e8e7513d78601a216d98eda95338bb60033456501135705014215498f330ef70033c5c601ae769357f5030605336af500de96b29633c5da009357050202155d8d2a9833460601ce7f935786012216d18f3386f601b38bc70033457501935605014215558d2a98b3c50701ee7793d6f5038605b3ead5003e9c769cb345890193d605028215d58dae98b3c41e01926613d68401a214458eb304dc0033099600b3c5250193d40501c215c58dae98334616019354f6030606458eea97b2973d8f935407020217458f3a9833460601935486012216458ee697330cf60033478701935407014217b36e97007698334606011357f6030606aa74598e7ae332f6da94ce94258d135605020215518d3306150133c7c900935787012217d98f33875400b389e70033453501935405014215b36895004696b2ea3d8e1355f6030606b367a6005e93529333c565009355050202154d8daa93b3457a0013d68501a215d18d3306d3003383c50033456500935605014215b362d500969333c575009355f5030605b366b500ca9fd69f3345ff01935505020215c98d2e9e33c5ca01ea74135685012215498e33859f00330fa600b3c5e50193d40501c215cd8c269eb345c6014a6613d5f5038605c98d62963e96b18c13d504028214458daa93b3c77700ae7413d78701a2175d8f26963a9632e6318d135605014215518d2ae31e95aaee398d1356f5032a670605518d2afa4e97369733c5ee00135605020215518d2a9e33c6c601ea669357860122165d8eba96b29636ea358d935605014215558daaf67295aaf2318d1356f5038e760605518d2afe9a96ae9633c5d800135605020215518d2a98b3c505010e6613d78501a215d98d36962e9632ee318d135605014215518daafa4295aae62d8d9355f50306054d8daae23275ca75aa95fa9533c6b200d666135706020216598eb296358d0a779357850122155d8dba95aa952ef2b18d13d60501c215d18daefeb695aeea2d8d9355f5030605c98da8022ef6a1451060833605fc1861358e398e10e0fd1521052104f5f5be701e74fe645e69be691e6afa7a5a7bba7b1a7cfa6c5a6dba6d7d618280197186fca2f8a6f4caf0ceecd2e8d6e4dae05efc62f866f46af06eec906103bc8500329c636fcc34aa8988699376f50093b616003337a000f98e6380063a814a89466368d5008d462a87850a0581e3ede6fe83cb85013285d68597000000e780a03b6365ac322a8d1305000463f5aa323305ac4133555501814c89456368b5008d452a86850c0581e3edc5fe938d2c0063ea9d316145b3b5ad02639a0530b384ad02ea9463eaa43113893c006a847d19268a630d0902630c0d24233044015285639b0b00130600105285814597400000e78060200860610408e1c10408e5e3f844fd17a5ffff13052506a5ac4ee0638b0d2e014b13098d0093891c005a85ee8597000000e780a03563030d201d05935435002330490163990b0052858145268697400000e780201bd29463e24425638669016109050b268ad1b7094963e72d0593098d02330a904105442285ee8597000000e780c0301d05135b350023b0990063990b00268581455a8697400000e780801633856401636195200504b3058a00e109aa84e39325fd11a02685d68597000000e7806028636fac2463860d262a8b938bfdff2a84638b0b161385edff9305f00363eda520854c5a846ae86ee463080d14aa843395ac00331d55013309a401636589186145b38da402c265ae9d3385ab022e9593098500130a0501636f2c0d03b50d000c612300b40013d68503a303c40013d605032303c40013d68502a302c40013d605022302c40013d68501a301c40013d605012301c400a181a300b40093558503a307b400935505032307b40093558502a306b400935505022306b40093558501a305b400935505012305b40093558500a304b4002304a4000c6180e500e15a85d6852686a28697000000e780c022058915ed5a85d6855e86a28697000000e780802183b5090013563500b295838605001d893395ac00c98e2380d50083350a00b29503860500518d2380a5004a846a99e37489f249a82685a26597000000e780c0185a85d6852686a28697000000e780801c83b58d0013563500b295038605001d893395ac00518d2380a50081cc1385f4ffa68b426de31c0dea97200000e78020b00000426da26d63638c0a33058c40826523b0650123b4850188e923bca50123b0b50323b45503e6704674a6740679e669466aa66a066be27b427ca27c027de26d0961828017a5ffff1305a5def14597200000e780e08e000017a5ffff130565ddf5b717a5ffff1305c5dccdb717a5ffff130525dce1bf17a5ffff130585d5ada817a5ffff1305e5d793054002c9b717a5ffff130505da5dbf17a5ffff130565d0a1a817a5ffff1305c5d84db717a5ffff130525d291a017a5ffff130585cb9305300271b717a5ffff1305a5da29a85285d68597000000e780c002637bac0017a5ffff130585dd97000000e7804005000017a5ffff1305e5cd9305100289bf01cd1306000463f0c5027d153355b50005053315b500828017a5ffff130585cb9305100239a017a5ffff1305a5cd9305400297200000e780c080000097200000e780e09c000063efa5006382a5021345f5ffaa951305000463f2a50205453315b500828017a5ffff1305c5c629a017a5ffff130525c69305100239a017a5ffff130545bf9305300297100000e780607b000063e0a6041307f003636cc7001307000463fde500898e33d5c6003355b500828017a5ffff1305e5c429a017a5ffff130545c49305400297100000e7806077000017a5ffff130565cfb545f5b790659461137806fc3698636bd80c98699355660063e3e500ba8594e2094694e6b68763ebc508fd1593d8860393d2060313d3860293d3060213de860193de060113df8600b68736863e879387070463efe7062380c70013578603a383e700135706032383e70013578602a382e700135706022382e70013578601a381e700135706012381e7002182a380c7002384d700a387170123875700a386670023867700a385c7012385d701a384e70190621ce6fd159ce23e86c9f99385070463e7f50214e1233405010ce914ed828017a5ffff130565b8f14597100000e780a068000017a5ffff130525b7f5b717a5ffff130585b6cdb7717106f522f126ed4ae94ee552e1d6fcdaf8def4e2f0e6eceae82a841305000497550000138ae5436371850417550000930425438860631e05348864fd558ce063130512c870cc6cd068d464aae4aee032fc36f80a850c1897000000e780209c054588e413850401c5a803350a04631b053203358a04fd552330ba041ded03350a0883358a0703360a07aae02efc32f80a850c1897000000e78080e705452334aa040265a2654266e2662338aa04233cba042330ca062334da0603398a0663000902033509000c6110650ce20c6510610ce6130b0a04630825032a8991a403390a0603358a056373a902130509046368252983350a042330aa0685052330ba046315092209a823340a0619ac03350a0405052330aa0403350a00631e052803358a00fd552330ba001ded03350a0a83358a0903360a0983368a08aae4aee032fc36f80a850c1897000000e780408d05452334aa0013050a018a851306000397400000e780c0c583398a031305f003636335210545814c3315350163788500850c63840c1c0605e36c85fe83350a0363e3bc00e68503358a020146e146b386dc02aa96138406fdb385bc406389c516630d051c147803b9060061047d16e307d9fe033509008335890088e1033589008335090088e5047017550000130b852803350b0183358b03934af6ffe69a5686ca8697000000e78000cd93553500a695038605001d89854b3395ab00518d2380a50063f85c11130c000417550000130b6524138afaff63778a1333954b01b3143501ca9463e72413033d840203350b0183358b035686ca8697000000e780a0c793553500ea95038605001d893395ab00518d2380a500833a840003350b0183358b035286ca8697000000e780c0c493553500d695038605001d893395ab00518d2380a50008600c612380b40013d68503a383c40013d605032383c40013d68502a382c40013d605022382c40013d68501a381c40013d605012381c400a181a380b40093558503a387b400935505032387b40093558502a386b400935505022386b40093558501a385b400935505012385b40093558500a384b4002384a4000c6184e504e12114d28ae3e54cf119a00149528b03350b0005052330ab004a85aa700a74ea644a69aa690a6ae67a467ba67b067ce66c466d4d61828017a5ffff1305658121a81795ffff1305c5749305300231a01795ffff1305e57ff14597100000e780203000001795ffff1305a572f9bf1795ffff1305057ecdb797100000e780204a000017a5ffff1305d5b49795ffff9386c56d15a017a5ffff1305b5b39795ffff9386a56c09a817a5ffff130595b29795ffff9386856bc1450a8697100000e78020450000317106fd22f926f54af14eed52e956e55ae1defce2f8e6f4eaf0eeec97550000938ce50683b50c04639d05382a8903b58c04fd5523b0bc041de9175500001304050548602c7c3078aae4aee032fc28002c1897000000e78060ae054528e42265c2656266827628e82cec30f034f403b50c0583b58c053335a9001345f5ffb335b9006d8d51c517550000130545002c75638e052090612300c90093568603a303d900935606032303d90093568602a302d900935606022302d90093568601a301d900935606012301d9002182a300c90013d68503a307c90013d605032307c90013d68502a306c90013d605022306c90013d68501a305c90013d605012305c90013d68500a304c9002304b900906165a203b50c0483b50c00050523b0ac04639b052a03b58c00fd5523b0bc0015ed175500001304c5f548704c6c50685464aae8aee4b2e036fc28002c1897f0ffffe780c04f054508e4130504012c001306000397400000e780608883ba0c03638f0a2283b98c02138afaff13848902854463809a04638b0922033b040003b50c0183b58c032686ca8697000000e780609593553500da9583c505001d8933d5a50005898504610469d5f91463e6440139a263030a108144930a0004268b63e49a00130b000483bb8c0303bc0c0161453385a4024e9513048502054d03b50c0183b58c032686ca8697000000e780808f638e091a833504fe13563500b2950386050093767500b316dd0093c6f6ff758e2380c500937515003306b040833604fe13661600329513563500369603460600937675003356d600058a51e2630b9b1263fe5b1333159500331575016295636e85131061146590e21065146190e691c12a89833d040003b50c0183b58c0385042686ca8697000000e780c08693553500ee95038605001d893315ad001345f5ff718d2380a5006104e3129af4d28405a023302901930585064a862334260123b02501930c050451a8638a090e814461453385a4024e9508610c612300b90013d68503a303c90013d605032303c90013d68502a302c90013d605022302c90013d68501a301c90013d605012301c900a181a300b90093558503a307b900935505032307b90093558502a306b900935505022306b90093558501a305b900935505012305b90093558500a304b9002304a9000c6123b425012330250103b50c00050523b0ac00ea704a74aa740a79ea694a6aaa6a0a6be67b467ca67c067de66d296182801795ffff1305c53429a01795ffff130525349305300231a01795ffff1305453ff14597100000e78080ef00001795ffff1305053893051002edb797100000e780e00900001795ffff130595749795ffff9386852d09a81795ffff130575739795ffff9386652cc145300097100000e780000600005d7186e4a2e026fc4af84ef452f056ec83ba050263800a0a2e8a2a898065b35954034e8597000000e780200b83340a002ae02ee402e863e335078145636e54031396350032950d466370560983c6140003c70400a206d98e03c7240083c7340033045441d6944207e2075d8fd98e14e185052105e37a54fd2ee8226502662338b9002334a9002330c900a6600664e2744279a279027ae26a616182800a8581454e8697000000e7806008c2650265e37954f9d9b71795ffff13054539e54597100000e78080de00001145d68597100000e780e0570000011106ec22e826e42a841dc51355c40305ed93351500931434008e0599c4268597200000e780800eaa8581e9268597200000e780a00f0000a1452e85a285e2604264a2640561828097d0ffffe780401b0000411106e497000000e78000037d567e1605066315c500a2604101828011e597d0ffffe780c01800002e8597200000e780c00a00005d7186e4a2e026fcae86b29563f4d5000145a1a82a8408659314150063e39500ae84914563e39500914493d5c40393b51500139634008e0501c914600e0536f0a14636f42af811a002f42800141097100000e780606aa265426599c1e26531a008e004e47d557e150505a6600664e27461618280411106e4054697000000e78060f87d567e1605066315c500a2604101828011e597d0ffffe780200e00002e8597200000e78020000000797106f422f026ec4ae84ee452e06365d7046366e604aa89b304d7403389d5002685814597100000e780806b2a842e8aca85268697300000e780a03b23b0890023b4490123b89900a2700274e2644269a269026a456182803685ba8519a03a85b28597100000e780203e0000797106f422f026ec4ae84ee452e06363d604aa89b304d6403389d5002685814597100000e78000652a842e8aca85268697300000e780203523b0890023b4490123b89900a2700274e2644269a269026a456182803685b28597100000e7800038000063e8c60063e9d500b385c640329582803285b68511a0368597100000e780e0350000011106ec22e826e42a8410690865ae846319a6002285b28597000000e78020ec10680860931536002e9504e1050610e8e2604264a26405618280397106fc22f826f44af04eec52e856e4114a32892a84637d46032d45ad4a814597100000e7802059aa84ae891795ffff9305e5132d46268597300000e780c028054508c0233444012338240104ecb1a803c5150003c6050083c6250083c535002205518dc206e205d58db3e4a500b9c09104638424052d45ad4a814597100000e78060532a8aae891795ffff9305250e2d46528597300000e78000232320040004e423382401233c4401233034032334540331a0114a631d4901154508c0e2704274a2740279e269426aa26a216182802d45ad4a814597100000e780c04daa84ae891795ffff930585082d46268597300000e780601d23200400a9b71061833805011c65210605483e8763ee17019307f7ff10e11ce5637d1801833686ff0c622106e3f3d5fe333517011345150082800545854597100000e780601e0000411106e410610e069796ffff938626d2369610620286907588711c6e9795ffff9385950d3d4635a8907588711c6e9795ffff9385c50b2d462da021052ae01795ffff9307c5071795ffff130745083d463da0907588711c6e9795ffff9385a5042146a2604101828721052ae01795ffff9307c5001795ffff1307e5001d468a862e85be8597100000e780000ca2604101828082808365050005466345b60099c9054609a809466389c5000d466394c500210521a0610511a041050c6591c5086117230000670083cb8280397106fc22f83287ae862a8402f002ec02e802e4130500022af405659b0815822c108d472800894201460148730000006309550285456308b502914515e522751306000289456361a602130514002c001306000297300000e78080062300040009a8854511a081450ce408e805452300a400e270427421618280397106fc22f83287ae862a8402f002ec02e802e4130500022af405659b0815822c109547280089420146014873000000630b55028545630cb502914515e922751306000289456365a602130524002c001306000297300000e780e0fe01458545a300b40009a80145a300040029a081450ce408e805452300a400e270427421618280130101ba233c1144233881442334914423302145233c3143233841432334514323306143233c7141b289ae8b2a8408081306004093040040814597300000e78080eb2338914005659b08c58293050141080889440146de864e8781470148730000006301950885456300b508914535ed03390141130500406372250b8545054b4a8597100000e780c0222a8aae8a0c081306004097300000e780c0f2930209c013050a402338514085659b88c58293050141130600408944de864e87814701487300000063019508630e6507114b25ed03350141094b63e8a2062330440123345401b1a8854511a081450ce408e8233004008330814503340145833481440339014483398143033a0143833a8142033b0142833b81411301014682804a85814597100000e780e018aa84ae890c084a8697300000e78000e904e0233434012338240145bf014b2334640108e823300400e3810afa528597200000e780c0a551bf9308d0057d558145014681460147814701487300000001a0086101a08280797106f42e8813564500130f7002130710279796ffff938e26e16363e608130f700213076102174600008338064939661b03068f05669b03b6479302c0f937e6f5051b0ef60faa86333515032d813b066502b307d600139607034992330676029355160141821376e67fbb855502be95769683471600c615c19103460600a30ff7fef69583c7150083c50500711f230fc7fea300f7002300b7007117e365defa130630066370a60493150503c99105661b06b647b385c502c5811306c0f93b86c502329546154191791f7695034615000345050093061100fa96a380c6002380a6002e85a945637cb5009305ffff130611002e961b0505032300a60005a006059305efff7695034615000345050093061100ae96a380c6002380a60093061100ae96130770020d8f1795ffff9305e50b4285014697000000e780e000a27045618280597186f4a2f0a6eccae8cee4d2e056fc5af85ef462f066ec6ae86ee4aa8403654503ba893689328aae8b937c1500b70a110063840c00930ab00293754500ce9c89e5814b8c6085e5a1a08145630e0a005286de86038706008506132707fc134717007d16ba957df6ae9c8c6095c103bd840063ffac01218925ed83c58403054633059d41634cb60af9e1aa8c2e85c9a0807084742285a6855686de86528797000000e7806014054b0dc15a85a6700674e6644669a669066ae27a427ba27b027ce26c426da26d656182809c6c2285ca854e86a6700674e6644669a669066ae27a427ba27b027ce26c426da26d6561828780581305000383c584032ee003bc040283bd840288d8054b238c64036285ee855686de86528797000000e780e00c51f5228a33049d4105047d1451c803b60d02930500036285029665d985bf09466398c50093051500058193dc150011a0814c03bc040203bd84028458130415007d1409c803360d026285a68502966dd9054b2dbf37051100054be389a4f26285ea855686de86528797000000e780e00511fd83368d016285ca854e86829619f5b30990417d5a7d59338529016309450303360d026285a6850296050975d50da083b68d016285ca854e868296e31005ee014b23a844030265238ca402c1bd6689333b9901e1b5797106f422f026ec4ae84ee49b070600370811003a89b6842e84aa896389070114704e85b2858296aa85054591ed81cc1c6c4e85a6854a86a2700274e2644269a269456182870145a2700274e2644269a269456182805d7186e4a2e026fc4af84ef452f056ec5ae85ee483320500146933e7d2003289ae896304072a638706101c6d8146338e29018507370311009308f00d1308000f4e8601a893051600918eae962e866303640efd17adc7630fc60d8305060013f4f50fe3d105fe834516009374f40113f7f50363fa8802834526001a0793f5f503b363b7006367040383453600f614ad909a0393f5f50333e4b300458c630c64089305460055b79305260013946400598c61bf93053600b20433e4930071b7630bc6078305060063d3050493f5f50f1307000e63ede5021307000f63e9e50203471600834726001377f70393f7f70303463600f615ad9132079a075d8f1376f603598ed18d370611006386c50285c263fd2601b385d90083850500130600fc63d7c500814591e539a0e39d26ffce8599c13689ae89638b021803388500930500026372b902814e63060916ca85ce86038606008506132606fc13461600fd15b29efdf581aa13877900619b3386e940b308c90093f678008145630d3701ce87038407008507132404fc934414000506a6957df6014691ce93f788ffba9783840700850793a404fc93c41400fd162696fdf693d638009747000083b7e7f89744000083b2e4f8b714001092048504939804018508b30eb6001da013173e001a97b386c34113763e00b3f45500a181b3f55500a695b3851503c191ae9e2deaddcab6833a839305000c368e63e4b600130e000c9375ce0f139435001a94dddd81451a8745df146393c4f6ff9d8099821067c58efd8eb6959346f6ff9d82046b1982558e7d8e93c6f4ff9d829980c58e046ffd8e3696b29513c6f4ff1d829980458e7d8e13070702b295e31d87fabdb7630803029305000c63e4b3009303000c814593f633008e06106021041347f6ff1d831982598e7d8ee116b295f5f611a0814533f65500a181b3f55500b295b3851503c191ae9e63fc0e01834685030546b305d8416345d60285ce814a25a80c7508719c6dce854a86a6600664e2744279a279027ae26a426ba26b6161828709466398c600138615008581935a160019a0ae8a8145033b0502833b85020459138415007d1409c803b60b025a85a68502966dd9054a81a037051100054a638ca40283b68b015a85ce854a86829605e533095041fd597d5433058900630a350103b60b025a85a6850296050475d511a05684333a54015285a6600664e2744279a279027ae26a426ba26b61618280411106e497000000e780801c0000197186fca2f8a6f4caf0ceecd2e8d6e4dae0b2891306000232f80d46230cc10203b4090202e002e82af02ef461c003b589026307051083b409009305f5ff8e058d8113891500a10493058003330ab5026104854a17050000130b458a906001caa276027583b584ff946e829665ed08482ad803058401230ca1024c4803b509012eda033684ff0c6001ce631756019205aa95906563046601014621a08c618c61054632e02ee4033684fe833504ff01ce631756019205aa95906563046601014621a08c618c61054632e82eec0c6492052e95106508618a85029649e5c104130a8afc13048403e31b0af6b1a003ba890163080a0483b4090103b409001305faff12051181130915002104a104120a106001caa2760275833584ff946e829639e1906003b584ff8a8502960ded4104411ac104e31e0afc03b589006368a9002da0014903b589006371a90203b5090012092a99a27602758335090003368900946e829619c1054511a00145e6704674a6740679e669466aa66a066b09618280907588711c6e9785ffff9385b5532d468287907588711c6e9785ffff9385455339468287411106e497000000e78080010000411106e497000000e780a0000000411106e497c0ffffe780401c0000757106e5014730012948bd4821a89306f6ff13d547009a92a30f56fe0507368663fcf800aa879372f50013030003e3e002ff13037005e1bf13050008198d130610086370c5021785ffff9307e55009462e85be8597000000e7800082aa60496182809305000897000000e78040560000757106e522e1a6fccaf8cef4d2f0d6ecdae8dee4e2e066fc6af86ef432892e8a014c814c81499745000003bba5b69745000083bba5b69745000083b4a5b600690c612ef008652aec13058a002ae01785ffff130525482ae8294d22e40da03305b6000345f5ff5915133515002300a4006265146d02758296ee8c6311051213f5f90f631b051063758901e9a8636c890d33058941b3058a014146637fc50063022c0d81463386d50003460600630da6098506e319d5fe75a013867500937686ff3386b640ad8e93b6160013371600d98ea1c20146930605ff02676297b387c5009c6313c4f7ffa58fda9733747401e18f8defb307c7009c6313c4f7ffa58fda9733747401e18f95e34106e3f9c6fc31a83387d500034707006307a7038506e319d6fe930605ffe3f9c6fa6304c5062264b386c50083c606006386a6010506e319c5fe05a0b286e296138c1600e3f026f5d29603c50600e31ba5f38149e28de28a39a04a8c8549e68dca8a63872c030345040001c96265146d11460275c265829611ed33869a41b3059a01e39a9aed0145f1bd4a8c2264f9b7014511a00545aa600a64e6744679a679067ae66a466ba66b066ce27c427da27d49618280411106e41b8605009306000802c26376d6002302b100054671a01bd6b50019ee13d665001366060c2302c10093f5f50393850508a302b1000946ada01bd6050115e613d6c5001366060e2302c10013964503699213060608a302c10093f5f503938505082303b1000d462da81396b50275921306060f2302c1001396e502699213060608a302c100139645036992130606082303c10093f5f50393850508a303b10011464c0097000000e780e0d9a26041018280397106fc907594712ae032f836f4886d906994658c612af032ec36e82ee41785ffff930525320a85300097000000e780a0b2e27021618280086117030000670063d5411106e408611b8605009306000802c26376d6002302b100054671a01bd6b50019ee13d665001366060c2302c10093f5f50393850508a302b1000946ada01bd6050115e613d6c5001366060e2302c10013964503699213060608a302c10093f5f503938505082303b1000d462da81396b50275921306060f2302c1001396e502699213060608a302c100139645036992130606082303c10093f5f50393850508a303b10011464c0097000000e78060caa26041018280397106fc90759471986d32f836f43af0906994658c61086132ec36e82ee42ae01785ffff930585220a85300097000000e78000a3e27021618280357106ed22e926e54ae1cefcd2f8d6f42a840345050109c5833a04008544d5a0b2892e89033a840003654a03833a04009375450091e93336500163880a021785ffff9305e50f35a063960a0483358a0203350a02946d9785ffff9385850e094682961dc5814a854469a81785ffff9305650d83368a0203350a02946e05068296854441e103b689014a85d28502968da803254a038544a303910283350a0203368a022ee432e8930571022eec83250a0303068a0383360a0003378a0083370a0103388a01aaceaecc2300c10636f43af83efcc2e02800aae403b689011785ffff13052502aae82c104a85029619e9c6652665946d9785ffff9385650409468296aa8423089400850a233054012285ea604a64aa640a69e679467aa67a0d618280397106fc22f826f44af02a841c7508719c6f3a89b684829722e8230ca10002e4a30c01002800a6854a8697000000e78060eb22658345810139c50544b9e5834591017d1513351500c264b335b0006d8d05c103c54403118901ed8c748870946d9785ffff938515fc05460544829611ed8c748870946d9785ffff9385a5f4054682962a8419a03334b0002285e2704274a274027921618280411106e497000000e78040a200001785ffff9306850709462e85b68517f3ffff6700834c397106fc22f826f42e848c752ae40870946d9785ffff938585074546829622ec2300a10202e8a30001021785ffff1306050408082c0097000000e780e0de42658345010239c50544b9e5834511027d1513351500e264b335b0006d8d05c103c54403118901ed8c748870946d9785ffff938595ef05460544829611ed8c748870946d9785ffff938525e8054682962a8419a03334b0002285e2704274a27421618280757106e5014730012948bd4821a89306f6ff13d547009a92a30f56fe0507368663fcf800aa879372f50013030003e3e002ff13037003e1bf13050008198d130610086370c5021785ffff9307e5e709462e85be8597f0ffffe7800019aa60496182809305000897000000e78040ed0000797106f422f026ec4ae84ee42a8404690865ae893309b640058d6363250308602695ce854a8697200000e780e0e4ca9404e8a2700274e2644269a269456182802285a6854a8697000000e780c0000468f9b75d7186e4a2e026fc2e966368b6042a8408659314150063639600b284a14563e39500a14493c5f4fffd9119c5106032f0054632f42af811a002f428001410268697000000e780e003a265426581cdfd55fe158505630ab50009ed97c0ffffe78060aa000008e004e4a6600664e27461618280626597100000e780809b0000011106ec22e826e44ae03289aa8499cd2e84886605c18c6a91cd88624a8697100000e780009805e180e419a023b40400854521a8630409024a85a28597100000e780209575d1814588e423b824018ce0e2604264a264026905618280228565f5e1b703e6450308619376060189ea1376060219ea086117f3ffff6700c3ee086117f3ffff6700037b086117030000670063e3411106e422e02a8411c96347040289c9228597100000e780209009a8054501a88545228597100000e780808d19c9a285a26002644101828097c0ffffe780809b0000228597100000e780808d0000797106f422f026ec4ae84ee42a8904690865058d2e84636fb50283390900894533859900636cb4007d148145228697200000e78080bca2943385990023000500850423389900a2700274e2644269a269456182804a85a685228697000000e780e0008334090155bf5d7186e4a2e026fc2e966368b6042a8408659314150063639600b284a14563e39500a14493c5f4fffd9119c5106032f0054632f42af811a002f428001410268697000000e780e003a265426581cdfd55fe158505630ab50009ed97c0ffffe780008e000008e004e4a6600664e27461618280626597000000e780207f0000011106ec22e826e43284aa8499cd88660dc18c6a99cd8862228697000000e780e07b19ed85458ce431a823b40400854511a88545228597000000e78020797dd1814588e480e88ce0e2604264a26405618280411106e422e02a8408617d1508e005e90c70086c8c6182950870086511c5086c97000000e780e075087811c5087497000000e780007508647d1508e409c5a2600264410182802285a2600264410117030000670003735d7186e4a2e026fc4af84ef452f056ec83ba0501368a3289aa8963e3da00d28a806108687de1286c7d5610e8637c55010870106c98651c6d4e85b2854a86d286829761a08465306463edc400b386540163ee96082c683307b600636ec7086376d70208700c6c1074147c1c6d0a85268782970345010069e9a26563e8550f286c2ce824e426866367b50eb3b6c400918c33359500558d49e5338554016363950463e7a5080c7c63eca508b3059540639745090c74a6954a85528697200000e780c0a723b45901238009000868050508e8a6600664e2744279a279027ae26a616182801785ffff130585c311a81785ffff1305e5c229a01785ffff130545c2f14597f0ffffe780802e00001785ffff130515b59785ffff938605b6c1450a8689a01785ffff130505c69305f002d1bf1785ffff130515c893052003d9b7528597000000e780e0a400001785ffff130525d99785ffff9386a5ba9305b0021306710197f0ffffe780804300001785ffff1305c5bc71b71785ffff1305e5bd9305e00241b7034505000e051786ffff1306a6e12a969786ffff938606e6369598751062146188711c6fb6858287411110650c69b29563edc50008611069fd568582637dd60028616369b502410182801785ffff13056589a14535a01785ffff1305a5ab9785ffff9386a5ace145300097f0ffffe780c03a00001785ffff1305b5be9305600297f0ffffe780601e0000797106f422f0aa8502c2280050009146114497000000e78020de0345810011e942656319850203654100a2700274456182801785ffff1305c5c99785ffff938645ab9305b0021306f10197f0ffffe780203400001785ffff130575bab54597f0ffffe780e0170000797106f422f09c6185079ce19dc7b2962ee463e6c6022a8436e83aec280097000000e78080f16265c265226608e80ce410e0a270027445618280000000001785ffff130585a19305b00297f0ffffe780a0120000197186fca2f8a6f4caf0ceecd2e8d6e4dae05efc03bb050003370b00846594692a89130517002330ab006dcd5ae409072330eb0065cbb28a36f85af02e8597000000e78060f09385440063ef950caa892ef4081097000000e78000ef8d4563faa50c09811304f5ff63fe8a02938b1a0013952b0026956364950c2af4081097000000e78060ec2a8a63998b0233854401636c950a2ae863f649051785ffff13058596f1a015452304a900233009005a8597000000e78020c3b1a08a0a33859a002105636895082af4081097000000e780a0e7b385440163e39508aa892ee863644509338549412aec280097000000e78080df6265c26522662338a9002334b9002330c9005a8597000000e780c0bde6704674a6740679e669466aa66a066be27b09618280000000001785ffff1305a58d3da81785ffff1305a5a1b9451da81785ffff1305458c25a01785ffff1305a58b39a81785ffff1305058b11a81785ffff1305658a29a01785ffff1305c5899305b00297f0ffffe780e0fa0000397106fc22f826f42a8402e408083000a146a144a28597000000e78060ba0345010105e16265631f9502a264086097000000e78080b32685e2704274a274216182801785ffff130545a59785ffff9386c5869305b0021306710297f0ffffe780a00f00001785ffff1305a597b94597f0ffffe78060f30000397106fc22f826f42a84a307010008081306f10085468544a28597000000e780a0b2034501010de16265631095048304f100086097000000e780a0ab2685e2704274a274216182801785ffff1305659d9775ffff9386e57e9305b0021306710297f0ffffe780c00700001785ffff1305a590b54597f0ffffe78080eb00005d7186e4a2e026fc4af8ae842a898c69054632e002e402e889c90a8597000000e780c0910266426411a001442808a685a28697000000e78040a9034581011de5027563168504c2652266826688602338b9002334c9002330d900a6600664e27442796161170300006700c3a01785ffff130545939775ffff9386c5749305b0021306f10297f0ffffe780a0fd00001785ffff13055587c94597f0ffffe78060e10000011106ec22e826e49c692a84637df700b384e74063e3d400b684b306970063ede60263f7d7001545a300a400054531a8998e639dd4028c61ba953285268697100000e780c051014504e42300a400e2604264a264056182801775ffff1305656ef14597f0ffffe780a0da00002685b68597f0ffffe780005400005d7186e4a2e026fc4af84ef452f02e8483b905012a896145a14597000000e780000b59c1aa84086888e8086488e4086088e0054a52e402e802ec1314ba002800a28597f0ffffe780a07d13050006a14597000000e780a00731c923304501233445012338050004ed9775ffff938545790cf1a2650cf5c2650cf9e2650cfd23303505233405042338050420ed23340900233839012330a900a6600664e2744279a279027a61618280614519a01305000697000000e780a00300000c6591c508611703000067002301828017b3ffff6700630617b3ffff6700630617b3ffff6700630617b3ffff6700c30a97b0ffffe780200e00005d7186e4a2e026fc4af8ae84806590612a892800a28597e0ffffe78040390345810019c5426529e109452300a90029a805040dc09305910080e4130610024a8597100000e780c03aa6600664e2744279616182801775ffff1305c571f14597f0ffffe78000c4000097f0ffffe78020e00000357106ed22e926e54ae1cefcd2f8d6f4daf02e89aa8a2800d68597000000e78040f7034581008944630b951675cd0345210283451102034631028346410222054d8d4206e206558e518d83456102034651028346710203478102a205d18dc2066207d98ed58d82154d8daae40345a101834591010346b1018346c10122054d8d4206e206558e518d8345e1010346d1018346f10103470102a205d18dc2066207d98ed58d82154d8daae00345210183451101034631018346410122054d8d4206e206558e518d83456101034651018346710103478101a205d18dc2066207d98ed58d82154d8d2afc0345a100834591000346b1008346c10022054d8d4206e206558e518d8345e1000346d1008346f10003470101a205d18dc2066207d98ed58d82154d8d2af829a082e482e002fc02f803b58a010c6903b40a0113060002639bc5040c6108181306000297100000e78080650125854421e103b50a0210610818a28597e0ffffe7808025c279638f09120665627bc145637fb50263070b004e8597000000e780c0de8144130550032300a90011a08544050475c823b88a002685ea604a64aa640a69e679467aa67a067b0d6182804145814597f0ffffe780004b2a892e8a4146ce8597100000e780201b0345190083450900034629008346390022054d8d4206e206558e518d83455900034649008346690003477900a205d18dc2066207d98ed58d8215c98d03459900034689008346a9000347b9002205518dc2066207d98e0346d90033e7a6000345c9008346e90022068347f900498ec20603b58a02e207dd8e558e14651c610216598e3696be9533b7f5003a966304d6003337d60015ef0ce110e563070a004a8597000000e780c0cf63070b004e8597000000e780e0ce03b40a0131b71775ffff13052547f14597f0ffffe780609900001775ffff1305e545f5b71775ffff130545479775ffff9386c54b9305b002900897f0ffffe780c0b100000e059775ffff9385a5c72e950c6105458285094582800d4582801145828097f0ffffe78000b10000357106ed22e926e54ae1cefcd2f8d6f4daf02e8a2a8908100546814597e0ffffe780a002034501020dc12275c27597000000e780a0faea604a64aa640a69e679467aa67a067b0d61828003156102831541020356210283461102231ea104c205d18da274627503560104c27aaeccaae42318c104f5c603150105a6652314a1002ee013050002130b0002814597f0ffffe780a02e2a84ae89ac08194697100000e780a04313d58403a306a40013d504032306a40013d58402a305a40013d504022305a40013d58401a304a40013d504012304a40013d58400a303a4002303940013d58a03a30aa40013d50a03230aa40013d58a02a309a40013d50a022309a40013d58a01a308a40013d50a012308a40013d58a00a307a40023075401130564018a85294697100000e78040f68144631c6a01130600022285ca8597100000e78060379334150063870900228597000000e780e0b213057004e38f04ec0145e1bd3945d1bd130101c0233c113e2338813e2334913e2330213f233c313d2338413d2334513d2330613d233c713b93070002631df6503a8ab6892a8903c5950103c6850183c6a50103c7b5012205518dc2066207d98e558d03c6d50183c6c50103c7e50183c7f5012206558e4207e2075d8f598e0216518d2af003c5150103c6050183c6250103c735012205518dc2066207d98e558d03c6550183c6450103c7650183c775012206558e4207e2075d8f598e0216518d2aec03c5950003c6850083c6a50003c7b5002205518dc2066207d98e558d03c6d50083c6c50003c7e50083c7f5002206558e4207e2075d8f598e0216518d2ae803c5150003c6050083c6250003c735002205518dc2066207d98e558d03c6550083c6450003c7650083c575002206558e4207e205d98dd18d82154d8d2ae413050002854597000000e780a09d630505422a8413060002814597100000e780e0d01145854597000000e780a09b63080540aa84a301050023010500a30005002300050013050002930b0002814597f0ffffe78060092a8bae8a2c001306000297100000e78060d9228597000000e780e09713054a0063634537814597f0ffffe7808006aae2aee682ea2320412dd00588028c0597f0ffffe780e0ee338649018802ce8597f0ffffe780e0ed166ab6695664268597000000e7804093dae2d6e6deead2eecef2a2f68545130514032308b116636a8530814597f0ffffe780c000aae4aee882ec0d4597d0ffffe780007f2330a12c2334b12c2338012c99c1814511a8880597e0ffffe780e08c8335012d0335012c8e052e95c1450ce18335012dd6698505138409012338b12c6362342d0335812c6399a500880597e0ffffe78080898335012d033a012c13953500529500e19384150005042338912c630f04280335812c639ca4008805a68597e0ffffe78060868334012d033a012c939a340033055a0100e136752295636d85262ad47010a8002c1097f0ffffe780c0de033b812c7d556384a4026410a10a52850c61130485002ed4a8002c10268697f0ffffe78060dce11a2285e3930afe63070b00528597000000e78060819665801a33863501a80097f0ffffe780e0d913061117a800a28597f0ffffe780e0d8f66536762e96a80097f0ffffe780e0d7a669c66a3665666a11c5166597f0ffffe780007d167511c5766597f0ffffe780207c82e002fc02f802f40403c802801a1306c002814597100000e78060ae130680132685814597100000e78060ad1775ffff930515cb4146228597100000e78000b9370501011b0505022320a114233c012a88051306800f814597100000e78020aa88058c0297b0ffffe78000b6a8008c051306800f97100000e78040b5a800ce85528697b0ffffe780c0bd8802ac001306800f97100000e78060b3880513060004814597100000e78080a5033581229305000263eaa50a5a655de5033501229a653386a50032e3ba66b335b600b6952ee78345012399c1fd552eeffd55130610082eeb637dc5121306000800136309c500098e2295814597100000e78040a088028402a28597b0ffffe78060c321459305312c9060a38ec5fe93568600238fd5fe93560601a38fd5fe935686012380d50093560602a380d500935686022381d50093560603a381d50061922382c5007d15a104a1055dfd0336812228108c0597100000e780a0a62c10130600024a8597100000e780a0a563870a004e8597f0ffffe780e0638330813f0334013f8334813e0339013e8339813d033a013d833a813c033b013c833b813b1301014082801775ffff1305e58825a01775ffff1305458839a81775ffff1305a58711a81775ffff1305058729a01775ffff13056586f14597e0ffffe780a02900001775ffff130525d89775ffff9386a5da9305b002900297e0ffffe780a04200001305000211a0114597f0ffffe780005c00009305000897f0ffffe780e09f0000697106f622f226ee4aea4ee652e2d6fddaf9def5e2f1e6ed2e8a2a89014481490d45aae082e49304110501163335c00093b51500b36ab500130b1108894b7d5c88088c0097f0ffffe780e056034501056309751f6301051003c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8d2ae903c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8d2ae503c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8d2ae103c5140083c5040003c6240083c6340022054d8d4206e206558e518d83c5540003c6440083c6640003c77400a205d18dc2066207d98ed58d82154d8daafc63890a00dda002e902e502e182fc639e0a0ca81813060002d28597100000e780c0c5012579e1639a091628110d46a28597e0ffffe780e0852a7559c96a75ca752a76aae9aee5b2e1a8188c0197f0ffffe78020320305eb008305db000346cb00e6792303a10aa205d18d2312b10a03459b0083458b000346ab008306bb0022054d8d4206e206558e518d2ad103451b0083450b0003462b0083463b0022054d8d4206e20683455b00558e518d03464b00a20583466b0003477b00d18d834c0108c2066207d98ed58d82154d8d2aed11a081496a658a550316410a8306610a2af82edc231ec102230fd102630e8409050401b5638609060305e1038315c1036256c2762307a1022316b10232d436f0130511010c103d4697000000e78080734ee423089101a8182c00054697f0ffffe78060eb667535c92a658a656676aaf0aeecb2e8880897f0ffffe78080012334a9004e8597f0ffffe78000b7014531a01305a005a300a90005452300a900b2701274f2645269b269126aee7a4e7bae7b0e7cee6c556182801775ffff1305c5a4f14597e0ffffe78000f700001775ffff130585ac9305b002edb71775ffff1305a5a49765ffff9386a52f9305b002900897e0ffffe780200f0000717106f522f126ed2a8432e402ec02e802fc02f8a303010232f4aee02800aae40808aae813057102aaec28109305710297f0ffffe780c02d058901e9034571020dc9a300a40005450da888102c101306800397000000e7804063f954ca65881097f0ffffe780c02a058969d991ccfd14f5b7c26562660ce810ec2300a400aa700a74ea644d61828097a0ffffe780c02d00004d7186e6a2e226fe4afa4ef652f256ee5aea5ee662e2e6fdeaf9eef5b2842e8a2ae0014c814d8149814b1304110cfd5a3d4d32e82ee48801e285268697d0ffffe780c04f0345010c631e052863045c3103459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8d2ae90345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8d2ae503459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8d2ae10345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8daafca81813060002d28597100000e780c08c0125631305188801e285268697d0ffffe780004d0e6b630d0b1ece6c2e65637f9d15aaeceef04145814597e0ffffe7800076aa84ae8b4146da8597000000e780204683c5840083c9940003caa40083cdb40003c6c40003cdd40083c7e40083caf40003c3040003c7140003ce240083c6340003c8440083c3540083c8640083c2740063870b04268542f4c68496e01a896af01e8d52ec728a6ef8b68dcee4ba89b2e856fcbe8aae8b97f0ffffe78060fede85d687e27a46664e87a669ee86c27d528e626aea83027d4a838662a68822780675631f0514a20933e5b900420ae20db3e54d014d8d220db365cd0013960701e20a33e6ca00d18d821533e9a500131587003365650093150e0113968601d18d4d8d93958300b3e505011396080193968201558ed18d82154d8daaf093840cff130a0b012685814597e0ffffe7802065aa8cae8bd285268697000000e7804035e6e1dee5a6e928118c0197f0ffffe78020e60c1988618c65814baa7daaf4aef88549c264226afd5a3d4d666511c55a8597f0ffffe780e0f0050c91bb2e6586765de533e5790111cd638c0d024675a675026608f20cee14e2233426012338b6013da01305500382652380a50023b80500638f0d006e8597e0ffffe780a07401a81305200382652380a50023b80500b6601664f2745279b279127af26a526bb26b126cee7c4e7dae7d716182801765ffff13054562f14597e0ffffe78080b400001765ffff130505639765ffff938685679305b002301197e0ffffe78080cd00001765ffff1305b56a93059002e9b797e0ffffe780c0cd0000757106e522e1a6fccaf8cef4d2f02a89814432e402e81304910181153335b00093351900b369b500094a28082c0097f0ffffe780a0e30345810165d9630c451303459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8daaec0345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8daae803459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8daae40345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8daae0e39909ee880013060002ca8597000000e78080530125e31e05ec93f4f40f850413f5f40fe30795ec1765ffff13058547f14597e0ffffe780c09900002685aa600a64e6744679a679067a4961828071c693f7f50f2300f5003307c500a30ff7fe894663fcc60aa300f5002301f500230ff7fea30ef7fe994663f1c60aa301f500230ef7fea14663fac60893f5f50f9b9785003307a0400d8bad9f198e9b950701ad9f2a97719a1cc3b305c70023aef5fe63f5c6065cc31cc723aaf5fe23acf5fee14663fcc604137847005cc71ccb5ccb1ccf6108939807029396070293d8080223a2f5fe23a4f5fe23a6f5fe23a8f5fe33060641fd474297c69663f0c7020116937706fe93870702ba9714e314e714eb14ef13070702e31af7fe8280397122fc26f84af44ef052ec56e85ae45ee093f735006387074069c2aa8719a06303062a83c60500850513f735002380d7007d1685076df793f637003e87cdea3d48637dc804930806ff6378180133e8b700137878006304083093d84800138f1800120f2e9f2e87be86832e0700032e4700032387000328c70023a0d60123a2c60123a4660023a606014107c106e31eeffc85089208c695c6973d8a137886001377460093762600058a630c080083a8050003a84500a107a10523ac17ff23ae07ff11c798419107910523aee7fe6391061e09c603c705002380e7006274c27422798279626ac26a226b826b216182807d476379c70a094883c805009841638806290d486386061d9306c6fe03c3150003c8250093f306ff13843700938435009382330123801701a38067002381070113d94600ae92a687a28803a8170083a5570083a697001b53870103a7d7009b1f88001b9f85009b9e86001b5888019bd585019bd686011b1e87003363f3013368e801b3e5d501b3e6c60123a0680023a2080123a4b80023a6d800c107c108e39657fa9307190092073516b385f40033067640a29793780601137886009376460013772600058a6384080883cb050003cb150083ca250003ca350083c9450003c9550083c4650003c4750083c3850083c2950083cfa50003cfb50083cec50003ced50003c3e50083c8f50023807701a380670123815701a381470123823701a382270123839700a383870023847700a38457002385f701a385e7012386d701a386c70123876700a3871701c105c1076304080483c2050083cf150003cf250083ce350003ce450003c3550083c8650003c8750023805700a380f7012381e701a381d7012382c701a382670023831701a3830701a105a1079dc203c3050083c8150003c8250083c6350023806700a380170123810701a381d70091059107e30307e283c6050003c715008907238fd7fea38fe7fe890539b513f73700e31d07ec39b59306c6fe93f306ff1384170093841500938213012380170113d94600ae92a687a28803a8370083a5770083a6b7001b53870003a7f7009b1f88011b9f85019b9e86011b5888009bd585009bd686001b1e87013363f3013368e801b3e5d501b3e6c60123a0680023a2080123a4b80023a6d800c107c108e39657fa9307190092073d16b385f40033067640a297a1b593d84800938e18002e88033e88000333080085062334c7012330670041084107e3e5d6ff85089208c695c6973d8a01bb9306c6fe03c8150093f306ff13842700938425009382230123801701a380070113d94600ae92a687a28803a8270083a5670083a6a7001b53070103a7e7009b1f08011b9f05019b9e06011b5808019bd505019bd606011b1e07013363f3013368e801b3e5d501b3e6c60123a0680023a2080123a4b80023a6d800c107c108e39657fa9307190092073916b385f40033067640a29749b3aa8709b919ca0347050083c705007d166317f700050585057df6014582800345050083c705001d9d8280aa862e87b287630db50cb388c5403308c040b388a84006082e832a8e6372181b3346b5001d8a637fb50a63010612cdcb1386f7ff9d4563f8c51813061700b305c54093b5750093c5150093f5f50f638a0516b365e5009d896395051693f587ffba95033603002103210e233ccefee39a65fe13f687ff13f57700aa87b385c600329739cd0345070005462380a5006389c704034517000946a380a5006382c704034527000d462381a500638bc702034537001146a381a5006384c7020345470015462382a500638dc700034557001946a382a5006386c700834767002383f5003685828029ea3306f5001d8a65ca1386f7fffdd7b307c5007d5821a07d16e30106ffb305c70003c5050093f57700fd17a380a700e5f59d4763fac70ab2871d48e117b305f7008861b385f60088e1e369f8fe93777600cdd7fd173306f700834506003386f6002300b600f5b71376750041ca9385f7ffc9d72a867d5821a0fd15e38005f903450700050693777600a30fa6fe0507edf79d4763fcb704938885ff93f888ffa10833051601ba8703b807002106a107233c06ffe31aa6fe469793f77500130617008ddfba9711a005060347f6ff0505a30fe5fee31af6fe36858280cdba3685d5b713061700f9bfb287a5b73285ae8713061700e1f919b73e8625bf2a86be8549bfd182e6ad7f520e5108c9bcf367e6096a1f6c3e2b8c68059b3ba7ca8485ae67bb6bbd41fbabd9831f2bf894fe72f36e3c79217e1319cde05bf1361d5f3af54fa54b598638d6c56d340101010101010101ff00ff00ff00ff00fffefefefefefefe80808080808080800a0a0a0a0a0a0a0a0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000018cd0900000000000010000000000000040000000000000018bd01000000000000100800000000004000000000000000010000000000000060090100000000000000000000000000011101250e1305030e10171b0eb44219110155170000023901030e0000032e001101120640186e0e030e3a0b3b053f198701190000042e00110112064018030e3a0b3b05360b3f198701190000052e006e0e030e3a0b3b05200b0000062e001101120640186e0e030e3a0b3b050000072e006e0e030e3a0b3b0b200b0000082e011101120640186e0e030e3a0b3b0b360b0000091d00311311011206580b590b570b00000a1d0031135517580b590b570b00000b1d00311311011206580b5905570b00000c1d0031135517580b5905570b00000d2e006e0e030e3a0b3b0b3f19200b00000e2e011101120640186e0e030e3a0b3b0b3f1900000f1d0131135517580b590b570b0000101d01311311011206580b590b570b0000111d01311311011206580b5905570b0000121d0131135517580b5905570b0000132e006e0e030e3a0b3b053f19200b0000142e011101120640186e0e030e3a0b3b05360b3f190000152e011101120640186e0e030e3a0b3b053f190000162e0111011206401831130000172e0011011206401831130000182e001101120640186e0e030e3a0b3b0b0000192e011101120640186e0e030e3a0b3b0b00001a2e011101120640186e0e030e3a0b3b0500001b2e011101120640186e0e030e3a0b3b05360b3f1987011900001c2e001101120640186e0e030e3a0b3b0b3f1987011900001d2e006e0e030e3a0b3b0b870119200b00001e2e001101120640186e0e030e3a0b3b0b360b3f198701190000007000000004000000000008016f2900001c001143000000000000051200000000000000000000700e0000021e2d00000200000000039a420100000000000e0000000152c44b000078350000010b0200021e2d000002463c000004a8420100000000000e00000001521d0e0000028e010300000000c722000004000000000008016f2900001c00f915000088000000051200000000000000000000a00e000002da180000021f050000057d0c00002f16000002f90501067877010000000000020000000152f03200002b0c000002eb01025c3c000002ab30000005fa350000712300000593030105fa350000712300000593030105fa350000712300000593030105fa350000712300000593030105fa35000071230000059303010594280000c52100000593030105e52a00001946000005930301056b380000833700000593030105c50b0000f90300000536050105fa3500007123000005930301000002ad0c000002ab300000055f3f00007123000007010401055f3f00007123000007010401055f3f00007123000007010401055f3f00007123000007010401055f3f0000712300000701040105c43000002c17000007010401054d0b0000e934000007010401000005a6000000c14600000273040105d71200000841000002730401056c4500002b050000024905010506080000cc000000024905010505280000f9030000026106010002a7300000023512000002a431000007454800004e27000003d00100022c3e0000071013000010460000038e0107403b0000a730000003890107403b0000a73000000389010000029c48000002632e0000087a770100000000004201000001529b1500008a35000004d3030965000000ea770100000000000200000004f1360adc1800000000000004f1150972000000fc770100000000000200000004f2360ae91800004000000004f215097f00000044780100000000000200000004fd360af61800007000000004fd1509f300000052780100000000000200000004fd470b000100006c78010000000000020000000403011e0b8c0000007e7801000000000002000000040701360c03190000a0000000040701150b0d0100008c7801000000000002000000040701470b1a0100009a7801000000000006000000040f0133000002a30b000007412b0000713b000004430107be2d0000482900000443010002242900000ddb130000b11b000004870100023c4400000d0d470000ce380000042a010002501400000e4880010000000000700000000152032e0000a7300000049a0fd902000020090000049b1110521a00004e8001000000000008000000044e1d11bd1900004e800100000000000800000019f8020909410100004e80010000000000080000001bef5000000af70200005009000004511c09d01e000060800100000000000400000004511609090300006e80010000000000080000000451280f952100008009000004651412071b0000b0090000225901090af41a0000e0090000171209000000000002650700000d87320000b11b000004870100026f0700000ed8860100000000007000000001521f030000a7300000049a0fe5020000800d0000049b1110a61a0000de8601000000000008000000044e1d11bd190000de860100000000000800000019f802090941010000de86010000000000080000001bef5000000ae2030000b00d000004511c09dd1e0000f086010000000000040000000451160909030000fe86010000000000080000000451280fa2210000e00d000004651412131b0000100e0000225901090af41a0000400e0000171209000000000000021f4a000013370a00006c0a000008bd0601137f030000672e000008f606011311490000f44000000810070105b90c000023050000086e050114bc78010000000000e4010000015289020000e031000008de04030bbc040000da780100000000000c00000008e504130bc9040000f6780100000000000400000008ea04190bd6040000327901000000000002000000080a051a12e3040000d00000000817052411c31c00001a7a010000000000040000000880051211b01c00001a7a010000000000040000000ec702090bfc1e00001a7a010000000000020000000e6d020c000000127511000010010000081a051112d01c0000400100000894041212b01c0000700100000ec702090cfc1e0000a00100000e6d020c00000012ac1e0000d0010000080b05200b50010000ac7901000000000006000000139403160b6a010000c07901000000000004000000139503090012b91e000000020000080c05210b5d010000b27901000000000004000000139403160b77010000c47901000000000004000000139503090011e3040000de790100000000001a000000080e052411c31c0000e479010000000000040000000880051211b01c0000e479010000000000040000000ec702090bfc1e0000e479010000000000040000000e6d020c00000011681d000008790100000000001c00000008eb041610031d000008790100000000001c00000012310910f71c000008790100000000001c000000112009105b1c000008790100000000001c00000011874c10ce1b000008790100000000001c00000010533111011c000008790100000000001c0000000a940d0910311c000008790100000000001c0000000c321110c11b000008790100000000001c0000000f7c091220190000300200000ab0091d1062190000147901000000000002000000092b350927010000147901000000000002000000095352000012431c0000800200000ab1091510711c00001679010000000000080000000f541c10141d000016790100000000000800000010501609bf1d000016790100000000000800000011871f000009121c00002079010000000000020000000f54150000000000000000000015f67a010000000000780300000152c0470000f92d0000083c0512701f0000b0020000083e05170c631f0000e00200001483020f00111a1e0000247b0100000000000400000008470525110d1e0000247b010000000000040000001641033311d0190000247b0100000000000400000016080327116e190000247b0100000000000400000019e502090999000000247b010000000000040000001b62500000000011e81b0000287b010000000000da0000000847052311db1b0000287b0100000000006e0000000a8b010912861d0000100300000a5801100f741d000040030000128c190fcb1d000070030000122c1209201900004c7b010000000000040000000b260e09e31d0000647b010000000000040000000b321209ef1d0000707b0100000000000a0000000b391309fb1d0000867b0100000000000a0000000b412509d71d0000607b010000000000040000000b2e1000000011dd1c0000487b010000000000040000000a57011211b01c0000487b010000000000040000000ec702090bfc1e0000487b010000000000020000000e6d020c00000011861d0000b47b0100000000004e0000000a8c010910741d0000b47b0100000000004a000000128c1910cb1d0000b47b0100000000004a000000122c120920190000b47b010000000000040000000b260e09fb1d0000ec7b0100000000000c0000000b412509ef1d0000e07b010000000000040000000b391309e31d0000dc7b010000000000040000000b32120000000012331e0000a0030000084c051312581e0000d003000016b9010911271e0000027c010000000000120000001814010c10dd190000087c0100000000000400000016dc1f0bbe1a0000087c01000000000004000000195a010f000000000c7d1f000000040000084c051c11681d0000367c010000000000720100000859052310031d0000367c0100000000007201000012310910f71c00003c7c0100000000001e000000112009105b1c00003c7c0100000000001e00000011874c10ce1b00003c7c0100000000001e00000010533111011c00003c7c0100000000001e0000000a940d0910311c00003c7c0100000000001e0000000c321110c11b00003c7c0100000000001e0000000f7c091220190000300400000ab0091d1062190000487c01000000000002000000092b350927010000487c01000000000002000000095352000012431c0000800400000ab1091510711c00004a7c010000000000080000000f541c10141d00004a7c0100000000000800000010501609bf1d00004a7c0100000000000800000011871f000009121c0000547c010000000000020000000f54150000000000000010211d00005a7c0100000000004e01000011220910ea1900005a7c01000000000014000000113a270b840100005a7c0100000000000600000019d60d1f11041a0000607c0100000000000800000019da0d200bf7190000607c0100000000000800000019460617000b111a0000687c0100000000000600000019db0d240010f71c00006e7c0100000000001a000000114715105b1c00006e7c0100000000001a00000011874c10ce1b00006e7c0100000000001a00000010533111011c00006e7c0100000000001a0000000a940d0910311c00006e7c0100000000001a0000000c321110c11b00006e7c0100000000001a0000000f7c091220190000b00400000ab0091d1062190000787c01000000000002000000092b350927010000787c01000000000002000000095352000012431c0000000500000ab1091510711c00007a7c010000000000080000000f541c10141d00007a7c0100000000000800000010501609bf1d00007a7c0100000000000800000011871f000009121c0000847c010000000000020000000f54150000000000000010f71c00008a7c0100000000001c000000114735105b1c00008a7c0100000000001c00000011874c10ce1b00008a7c0100000000001c00000010533111011c00008a7c0100000000001c0000000a940d0910311c00008a7c0100000000001c0000000c321110c11b00008a7c0100000000001c0000000f7c091220190000300500000ab0091d1062190000967c01000000000002000000092b350927010000967c01000000000002000000095352000012431c0000800500000ab1091510711c0000987c010000000000080000000f541c10141d0000987c0100000000000800000010501609bf1d0000987c0100000000000800000011871f000009121c0000a27c010000000000020000000f541500000000000000102d1d0000dc7c01000000000012000000115a1209e91f0000e87c01000000000004000000117f0e0010ab1900000a7d01000000000006000000115019102b1a00000a7d010000000000060000001b1a0e117a1900000a7d0100000000000600000019e5020909a60000000a7d010000000000060000001b62500000000a2c190000b00500001150190a391d0000f005000011541b0f381900006006000011631a10861900007c7d01000000000002000000092b3509340100007c7d01000000000002000000095352000009451d00007e7d0100000000000c00000011641b10511d0000947d0100000000001200000011661609f61f0000a07d01000000000004000000117f0e00091e1a0000067d01000000000004000000114f2c1098190000f27c01000000000010000000114a12114b1f0000fe7c010000000000040000001bcb051b113d1f0000fe7c010000000000040000000d7e04080b2b1f0000fe7c010000000000040000000d2e030900000000000012e3040000b00600000863052811c31c0000047e010000000000040000000880051211b01c0000047e010000000000040000000ec702090bfc1e0000047e010000000000020000000e6d020c0000001175110000307e010000000000260000000865051512d01c0000f00600000894041212b01c0000200700000ec702090cfc1e0000500700000e6d020c000000000d3c380000ae2d000008f2011337170000372b000008f4050113263100001729000008430701051a270000431c0000089c0401167a850100000000009800000001526211000011f916000086850100000000001800000008e6071b0b6510000086850100000000000c0000001f1701120011c1160000ac850100000000005800000008e807091169210000b6850100000000004a0000001f65012711b5150000b885010000000000480000002027051611c9150000cc85010000000000060000001f66013c0bc9040000cc85010000000000060000001f700109000b65100000d485010000000000140000001f6701150b65100000ea85010000000000160000001f69011100000000131f0700005723000008e5070100021e1a000005f8160000fb2e0000089304010002012f000002e031000006a07a010000000000560000000152cf490000d819000008f304000005fa0800008b49000008640401051b0f00001f09000008790401157c7e0100000000007e010000015245390000fb2e00000838040c591000008007000008390419128b1c0000b0070000084d041d0a44190000e00700001d2f110012a9110000100800000856041a11b6110000047f01000000000018000000086b04150bb30100000a7f010000000000120000000881042c0011b61100002a7f01000000000018000000086c04190bb3010000307f010000000000120000000881042c0011381a00004a7f010000000000040000000873041f11ca1a00004a7f010000000000040000001996011a09b30000004a7f0100000000000400000017ee1c00000bbf0100004e7f010000000000080000000876040b0012971c000040080000083f041d0a50190000700800001d2f11000bcb0100009c7f0100000000000a0000000846041512451a0000a0080000085d042612d61a0000e0080000195a010f10e21a0000ca7f0100000000000400000017d93609c0000000ca7f0100000000000400000017ee1c0000000002f101000007d53c0000bd3800001f550102ec3700000eb880010000000000bc010000015292350000372b00001f1f0fab1d0000100a00001f201212981d0000400a0000123f050911971e00003e81010000000000d40000001272020f116c1a0000488101000000000008000000249e01320b251b0000488101000000000008000000195a010900116f1b00005081010000000000ac00000024a20122097b1b000056810100000000001a000000252c1010871b000070810100000000008c000000252f0510cd00000070810100000000000c0000002552160b8401000070810100000000000c0000000540051600109f1b0000b6810100000000000a000000256a160910200000b681010000000000020000002514070010931b0000a0810100000000000a0000002569160903200000a081010000000000020000002514070009da00000094810100000000000400000025651b097b1b0000e88101000000000014000000257716097b1b0000c88101000000000012000000255a1e000011791a000008820100000000000200000024b701430b251b0000088201000000000002000000195a010900111c1f00000a820100000000000400000024b8011c115c1b00000a82010000000000040000000da9050d093e1b00000a8201000000000004000000231a0900000000000f401e0000700a00001f252712841e0000a00a0000165f040d12711e0000d00a000024450229125f1a0000000b000024de0309110f1f00001a810100000000000a0000001909091311501b00001a810100000000000a0000000da9050d093e1b00001a810100000000000a000000231a09000000000000000002623d000002f644000005920400004e2700001f3501010002d119000005fc2200004e2700001f6501010000023d290000058f490000ae4600001f6f0101155a84010000000000200100000152bd090000f64400001f3401125c210000b00b00001f35012311a21500007e84010000000000de0000002027051612c9150000e00b00001f3601100cc9040000100c00001f700109000b65100000a684010000000000160000001f3801150c65100000400c00001f4101110b7c210000dc84010000000000020000001f41011112d4160000700c00001f3c01220f7f100000b00c00001f1a0911eb160000fc840100000000000a00000008a30412098a1f0000fc840100000000000a0000001f1a260000000b651000004885010000000000120000001f3e011100000013bd1c0000d11900001f6301010002b547000007821c0000b92d00001f15010002f108000002b92d0000071f3500004e2700001f1a0100000569310000ec2200001f1301010002e82f0000167482010000000000b400000001526b17000010b922000082820100000000009600000008a41a11a72200008282010000000000960000002679022a0c9a220000300b000026b6060f00000017288301000000000038000000015277170000074d180000ee2f000008a30107c5440000994b000008bf010002ab3000001860830100000000000a0000000152ef4700002842000008c6196a83010000000000b6000000015253420000ee2f000008ca106b1700007883010000000000a200000008cb0910b92200007a830100000000009600000008a41a11a72200007a83010000000000960000002679022a0c9a220000700b000026b6060f000000001920840100000000003a000000015296370000994b000008ce097717000040840100000000001400000008cf090000027809000005b40f0000a730000008bb09010002210c00001a20860100000000001600000001525f300000ff0f000008d0080b3d18000020860100000000001600000008d0083e000000028c39000002164a0000029548000019747701000000000004000000015282090000fd4b000001fa10a101000074770100000000000400000001fa05093400000074770100000000000200000003d21e0000000000029039000005f909000068100000065f0a0105f909000068100000065f0a0105f909000068100000065f0a0105f909000068100000065f0a010002b131000002fa1c00000279230000077a33000056450000097c0107c63a0000c1010000097c01076b2a000027410000097c0107b34a00000b3e0000097c0107f91a0000b73c0000097c0100024c3600000712000000fd190000094b01072b2d0000514900001b5b0107f5310000d52100001b5b0107e52100005f340000094b010002a94a00000503370000274100001bc705010002ab30000007c20a0000b03a00001b190100029b0b000007731b0000dd4100001bd901000002ab30000005641100002a1a000019e4020105a91a0000f62700001956010105f1430000e246000019cb0d010585250000ac3d00001998060105b3050000c33d0000194206010543410000b008000019860d010534280000802800001916040105f53700009f3a000019e402010553190000ab110000198f01010597410000432f000019560101051f2600002809000019f7020105a90d0000ca17000019040901054c040000a919000019560101054c040000a919000019560101020f0700000312860100000000000e0000000152ab4200007a390000190b0d00051f2600002809000019f702010002b403000002ec370000074a050000ed31000017d7010775340000f028000017e30107400d0000d911000017d70107353e00001231000017e30100028d37000005fa0100003646000017ec01010002ab30000007542f00006c17000017110107542f00006c1700001711010002623d000005c3140000ed310000175f0101000002ec0c00000259490000075a140000983b00002352010002ab30000007b71b0000573d000023190107b71b0000573d0000231901000002b22d000007d8170000b22d000025290107a63b0000de3b00002534010d74470000341c000025470107760f0000a93e000025130107760f0000a93e0000251301000002fa1c000002242d000002b029000002494300000538120000842300000aaa090105663c0000ad3f00000a8f0d01058f360000f60000000a560101053a080000ba0e00000a8a0101000002801000000286100000075a2700009b3900000c310102b50c00000780400000901000000c35010000000002b846000002712e000002ec37000007752e0000ff1c00000f78010002304a0000075e4300001c1f00000f5401000002294a000002ec370000077907000078120000104d01020c000000025f4500000744160000590000001050010000000002ef1a000002f108000007fe050000db2500001d2e0107461300002c2200001d2e01000000022d08000002ec3700000593450000ca2000000e6c02010002cc46000005db200000274100000ec6020105db200000274100000ec6020105db200000274100000ec602010000000208000000020c0000000d760a0000e519000011860107270e000052430000111a0102e519000007be1e00004e270000118701000d790800004419000011260107d03d0000fd120000117a0107242a0000d201000011720107242a0000d201000011720107d03d0000fd120000117a010002fa1c000002ab30000007a04800000c00000012300107394a00001f01000012290100025949000007331a00001f010000128a010002cf2f00000570260000b00b0000126c020100020b42000005e22b0000dd2f0000123e0501000002b60a0000076b3d0000a53c00000b180107b9290000d63600000b240107dc0e0000f82900000b0b010770210000b22100000b11010770210000b22100000b11010770210000b22100000b11010002ab3000000551360000f73300001607030105b0270000d54600001640030107f60c0000082a000016d30105fd3300003934000016b80101050a040000473d0000165b04010002242d000002bb300000052401000046050000181301010000025f4700000224290000052d4b00006747000024dd03010002cc46000005be26000067470000244102010002ab30000005642c00003a320000249b0101000000026845000005673a0000101a0000138f030105b73100005b0e0000138f0301027c2b00000244140000056e4400000347000021e80101056e4400000347000021e8010100000002ec0c000002f00c000002ec00000005df180000f43300000d5305010002e322000005d43800002e2900000da8050105d43800002e2900000da80501000005464400000a2f00000d930401027f3700000562490000192a00000d2a03010005cc080000192a00000d7d040100023308000002b4300000057d0e0000370500001456020105b4430000903a00001482020105ba0300003341000014bb03010591060000f50d000014120601001b2c800100000000000e00000001522c3f00006c390000148b070311492000002e800100000000000c000000148c0705093d2000002e800100000000000c0000001c8605000000029c480000023c44000005662d0000f64600001ae4040105662d0000f64600001ae4040105664600008c4b00001acd040105664600008c4b00001acd0401000002e62800001c6e7e0100000000000e0000000152cc150000fd2d00001c6e1d113d0000e31100001c95011d450f00005f3100001c85011e3a800100000000000e000000015224300000154200001c50030002a4190000021526000015fa7f010000000000120000000152fc440000a73000001ebb021172100000fa7f010000000000120000001ebc021b1137130000fa7f01000000000012000000084407090965100000fa7f010000000000120000001f5912000000000230320000150c80010000000000120000000152c2020000a73000001ed60211721000000c80010000000000120000001ed7021b11371300000c80010000000000120000000844070909651000000c80010000000000120000001f5912000000000002d4130000031e800100000000000e0000000152ec040000f711000020720602ae4700000545320000801800002025050105cd060000eb3b00002025050100021a30000005bc3e00005b090000209b07010000026a26000002c01700000563220000892b0000225801010563220000892b00002258010100021a3000000e3686010000000000a2000000015207100000a730000022830f62110000f00c000022830a12f9160000200d000008e6071b0c65100000500d00001f1701120011c116000074860100000000005800000008e8070911692100007e860100000000004a0000001f65012711b51500008086010000000000480000002027051611c91500009486010000000000060000001f66013c0bc90400009486010000000000060000001f700109000b651000009c86010000000000140000001f6701150b65100000b286010000000000160000001f69011100000000000000028c060000021735000005db2c0000091800002699060105121800000e2d000026b5060102ab300000054c150000b94400002677020100000000003c0000000200000000000800ffffffff9a420100000000000e00000000000000a8420100000000000e0000000000000000000000000000000000000000000000bc0100000200740000000800ffffffff74770100000000000400000000000000787701000000000002000000000000007a770100000000004201000000000000bc78010000000000e401000000000000a07a0100000000005600000000000000f67a01000000000078030000000000006e7e0100000000000e000000000000007c7e0100000000007e01000000000000fa7f01000000000012000000000000000c8001000000000012000000000000001e800100000000000e000000000000002c800100000000000e000000000000003a800100000000000e0000000000000048800100000000007000000000000000b880010000000000bc010000000000007482010000000000b4000000000000002883010000000000380000000000000060830100000000000a000000000000006a83010000000000b60000000000000020840100000000003a000000000000005a8401000000000020010000000000007a85010000000000980000000000000012860100000000000e00000000000000208601000000000016000000000000003686010000000000a200000000000000d886010000000000700000000000000000000000000000000000000000000000ec77010000000000f077010000000000f477010000000000fc7701000000000008780100000000000c7801000000000000000000000000000000000000000000fe7701000000000006780100000000000c780100000000001478010000000000000000000000000000000000000000004678010000000000527801000000000054780100000000005e780100000000000000000000000000000000000000000080780100000000008c780100000000008e7801000000000096780100000000000000000000000000000000000000000036790100000000003c7901000000000040790100000000004679010000000000fa790100000000002a7a010000000000000000000000000000000000000000005a7a0100000000007a7a0100000000009a7a010000000000a07a01000000000000000000000000000000000000000000627a0100000000006a7a0100000000009a7a010000000000a07a01000000000000000000000000000000000000000000627a0100000000006a7a0100000000009a7a010000000000a07a01000000000000000000000000000000000000000000627a0100000000006a7a0100000000009a7a010000000000a07a01000000000000000000000000000000000000000000ac79010000000000b279010000000000c079010000000000c47901000000000000000000000000000000000000000000b279010000000000b679010000000000c479010000000000c8790100000000000000000000000000000000000000000008790100000000000c79010000000000147901000000000016790100000000001e790100000000002079010000000000227901000000000024790100000000000000000000000000000000000000000016790100000000001e790100000000002079010000000000227901000000000000000000000000000000000000000000f87a0100000000000e7b010000000000107b010000000000187b01000000000000000000000000000000000000000000f87a0100000000000e7b010000000000107b010000000000187b010000000000000000000000000000000000000000003a7b010000000000447b0100000000004c7b010000000000967b010000000000000000000000000000000000000000003a7b0100000000003e7b0100000000004c7b010000000000927b010000000000000000000000000000000000000000003a7b0100000000003e7b0100000000004c7b010000000000927b01000000000000000000000000000000000000000000027c010000000000187c0100000000001e7c010000000000227c01000000000000000000000000000000000000000000027c010000000000187c0100000000001e7c010000000000227c010000000000000000000000000000000000000000001a7c0100000000001e7c010000000000247c010000000000267c010000000000000000000000000000000000000000003c7c010000000000407c010000000000487c0100000000004a7c010000000000527c010000000000547c010000000000567c0100000000005a7c010000000000000000000000000000000000000000004a7c010000000000527c010000000000547c010000000000567c010000000000000000000000000000000000000000006e7c010000000000727c010000000000787c0100000000007a7c010000000000827c010000000000847c010000000000867c010000000000887c010000000000000000000000000000000000000000007a7c010000000000827c010000000000847c010000000000867c010000000000000000000000000000000000000000008a7c0100000000008c7c010000000000967c010000000000987c010000000000a07c010000000000a27c010000000000a47c010000000000a67c01000000000000000000000000000000000000000000987c010000000000a07c010000000000a27c010000000000a47c01000000000000000000000000000000000000000000107d010000000000127d010000000000567d0100000000005a7d0100000000005c7d010000000000627d010000000000000000000000000000000000000000001a7d010000000000227d010000000000247d010000000000287d0100000000002a7d010000000000307d010000000000327d010000000000427d010000000000447d010000000000467d0100000000004a7d010000000000567d01000000000000000000000000000000000000000000627d0100000000007a7d0100000000007c7d0100000000007e7d0100000000008a7d0100000000008c7d0100000000008e7d010000000000927d01000000000000000000000000000000000000000000ac7d010000000000b27d010000000000b67d010000000000bc7d010000000000e27d010000000000147e01000000000000000000000000000000000000000000387e010000000000407e010000000000527e010000000000567e01000000000000000000000000000000000000000000387e010000000000407e010000000000527e010000000000567e01000000000000000000000000000000000000000000387e0100000000003c7e010000000000527e010000000000567e01000000000000000000000000000000000000000000947e0100000000009c7e010000000000a07e010000000000a87e01000000000000000000000000000000000000000000ae7e010000000000d87e010000000000587f010000000000687f01000000000000000000000000000000000000000000ae7e010000000000d87e010000000000587f010000000000687f01000000000000000000000000000000000000000000ea7e010000000000f87e010000000000fc7e010000000000567f010000000000000000000000000000000000000000006c7f0100000000008a7f010000000000a87f010000000000b27f010000000000000000000000000000000000000000006c7f0100000000008a7f010000000000a87f010000000000b27f01000000000000000000000000000000000000000000b67f010000000000bc7f010000000000c27f010000000000c67f010000000000ca7f010000000000ce7f01000000000000000000000000000000000000000000b67f010000000000bc7f010000000000c27f010000000000c67f010000000000ca7f010000000000ce7f010000000000000000000000000000000000000000004e80010000000000a480010000000000aa80010000000000b880010000000000000000000000000000000000000000005e80010000000000608001000000000076800100000000007a800100000000000000000000000000000000000000000084800100000000008e80010000000000aa80010000000000b8800100000000000000000000000000000000000000000084800100000000008e80010000000000aa80010000000000b8800100000000000000000000000000000000000000000084800100000000008e80010000000000aa80010000000000b88001000000000000000000000000000000000000000000fe8001000000000016810100000000003681010000000000128201000000000000000000000000000000000000000000fe8001000000000016810100000000003681010000000000128201000000000000000000000000000000000000000000168101000000000024810100000000004282010000000000468201000000000000000000000000000000000000000000168101000000000024810100000000004282010000000000468201000000000000000000000000000000000000000000168101000000000024810100000000004282010000000000468201000000000000000000000000000000000000000000168101000000000024810100000000004282010000000000468201000000000000000000000000000000000000000000828201000000000086820100000000008e820100000000009482010000000000b082010000000000b682010000000000000000000000000000000000000000007a830100000000007e8301000000000086830100000000008c83010000000000a883010000000000ae8301000000000000000000000000000000000000000000708401000000000072840100000000007e840100000000005c8501000000000000000000000000000000000000000000828401000000000086840100000000008a840100000000008e8401000000000000000000000000000000000000000000828401000000000086840100000000008a840100000000008e8401000000000000000000000000000000000000000000cc84010000000000d684010000000000d884010000000000dc8401000000000000000000000000000000000000000000ea84010000000000ee84010000000000f48401000000000032850100000000003685010000000000408501000000000000000000000000000000000000000000ea84010000000000ee84010000000000f48401000000000032850100000000003685010000000000408501000000000000000000000000000000000000000000408601000000000042860100000000004486010000000000cc8601000000000000000000000000000000000000000000408601000000000042860100000000004486010000000000608601000000000000000000000000000000000000000000408601000000000042860100000000004486010000000000548601000000000000000000000000000000000000000000de8601000000000034870100000000003a87010000000000488701000000000000000000000000000000000000000000ee86010000000000f08601000000000006870100000000000a870100000000000000000000000000000000000000000014870100000000001e870100000000003a8701000000000048870100000000000000000000000000000000000000000014870100000000001e870100000000003a8701000000000048870100000000000000000000000000000000000000000014870100000000001e870100000000003a870100000000004887010000000000000000000000000000000000000000009a42010000000000a842010000000000a842010000000000b642010000000000000000000000000000000000000000007477010000000000787701000000000078770100000000007a770100000000007a77010000000000bc78010000000000bc78010000000000a07a010000000000a07a010000000000f67a010000000000f67a0100000000006e7e0100000000006e7e0100000000007c7e0100000000007c7e010000000000fa7f010000000000fa7f0100000000000c800100000000000c800100000000001e800100000000001e800100000000002c800100000000002c800100000000003a800100000000003a8001000000000048800100000000004880010000000000b880010000000000b8800100000000007482010000000000748201000000000028830100000000002883010000000000608301000000000060830100000000006a830100000000006a83010000000000208401000000000020840100000000005a840100000000005a840100000000007a850100000000007a85010000000000128601000000000012860100000000002086010000000000208601000000000036860100000000003686010000000000d886010000000000d8860100000000004887010000000000000000000000000000000000000000007261775f7665630073747200636f756e74005f5a4e34636f726535736c6963653469746572313349746572244c542454244754243134706f73745f696e635f73746172743137683231633736663939343638653065646545007b636c6f7375726523307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e005f5a4e34636f726533707472347265616431376831626239643039646638396234373532450077726974653c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e007b696d706c2335347d00616476616e63655f62793c636f72653a3a7374723a3a697465723a3a43686172496e64696365733e006e657874005f5a4e34636f726533737472367472616974733131305f244c5424696d706c2475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c5424737472244754242475323024666f722475323024636f72652e2e6f70732e2e72616e67652e2e52616e6765546f244c54247573697a652447542424475424336765743137683633326532303137643665353735396645006e6578743c5b7573697a653b20345d3e00636f6e7461696e735f6e6f6e5f636f6e74696e756174696f6e5f62797465006275696c64657273005f5a4e3131305f244c5424636f72652e2e6f70732e2e72616e67652e2e52616e676546726f6d244c54247573697a6524475424247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c54242475356224542475356424244754242447542435696e6465783137686163396536316662616530626263376145005f5a4e34636f726533666d7439466f726d617474657231327061645f696e74656772616c3137686238656639343965396131613633346545005f5a4e36335f244c5424636f72652e2e63656c6c2e2e426f72726f774d75744572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683636336332373865383138373636393045005f5a4e34636f726533666d74336e756d35335f244c5424696d706c2475323024636f72652e2e666d742e2e55707065724865782475323024666f7224753230246936342447542433666d743137683464336136353331313038303933376445005f5a4e34636f726533666d7439466f726d617474657239616c7465726e617465313768333537326537646636323036356664374500696e646578005f5a4e34636f7265366f7074696f6e31354f7074696f6e244c5424542447542439756e777261705f6f72313768343165333439646137383638346138334500616c69676e5f6f66667365743c75383e005f5a4e34636f72653373747232315f244c5424696d706c24753230247374722447542439656e64735f776974683137683139626662313333653233336465306145005f5a4e34636f726535736c69636532395f244c5424696d706c2475323024247535622454247535642424475424336765743137683233646638653962656438656665346645005f5a4e34636f726533666d74386275696c64657273313044656275675475706c65356669656c6432385f24753762242475376224636c6f73757265247537642424753764243137686363643963626231656235626135633645005f5a4e34636f726536726573756c743133756e777261705f6661696c65643137683030653934303161326339653536633045007074720070616464696e670077726974653c636861723e0069735f736f6d653c7573697a653e00676574005f5a4e37355f244c54247573697a65247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c542424753562245424753564242447542424475424336765743137683362336666656535366439303731313345005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243873706c69745f61743137683461343239666364306233623563343945005f5a4e3131305f244c5424636f72652e2e697465722e2e61646170746572732e2e656e756d65726174652e2e456e756d6572617465244c54244924475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e65787431376831623734616564656639323065303665450063686172005f5a4e34636f7265366f7074696f6e31354f7074696f6e244c5424542447542436696e736572743137686265366237313331636461646331646245005f5a4e34636f726536726573756c743139526573756c74244c542454244324452447542438616e645f7468656e313768316532623263316238653933626561654500636f70795f66726f6d5f736c696365005f5a4e34636f726533666d7439466f726d6174746572323564656275675f7475706c655f6669656c64315f66696e6973683137683963326264643732306464613133376545007b696d706c2332397d007b696d706c2336357d005f5a4e3130385f244c5424636f72652e2e697465722e2e61646170746572732e2e66696c7465722e2e46696c746572244c5424492443245024475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722447542435636f756e743137683631323362313132363938303130326445005f5a4e34636f72653370747235777269746531376830336462313664353065636536366165450072616e6765006f7074696f6e005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f72336e74683137683635613666633036633265613031396645005f5a4e34636f72653373747235636f756e743134646f5f636f756e745f6368617273313768653066306166323562653730356463664500616c69676e5f746f5f6f6666736574733c75382c207573697a653e005f5a4e34636f726533636d70336d696e3137683961303232643031326665326338333745007b696d706c23317d005f5a4e34636f726533666d743372756e313768666639613633333362396633663061614500676574636f756e7400697465725f6d75743c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e006272616e63683c28292c20636f72653a3a666d743a3a4572726f723e007b696d706c2332357d005f5a4e34636f7265336f70733866756e6374696f6e36466e4f6e63653963616c6c5f6f6e63653137683331326365396462383432326365623645005f5a4e34636f726533666d74386275696c64657273313044656275675475706c65356669656c643137686134393061356537663734366534656245005f5a4e34636f72653130696e7472696e736963733139636f70795f6e6f6e6f7665726c617070696e673137683165326664363834393232323263326345005f5a4e34636f726533666d7439466f726d6174746572397369676e5f706c75733137683765363563323535316433616561343445007369676e5f706c7573005f5a4e34636f72653373747235636f756e743233636861725f636f756e745f67656e6572616c5f6361736531376864313333363866323830386530613030450076616c69646174696f6e73005f5a4e34636f726535736c696365346974657238375f244c5424696d706c2475323024636f72652e2e697465722e2e7472616974732e2e636f6c6c6563742e2e496e746f4974657261746f722475323024666f7224753230242452462424753562245424753564242447542439696e746f5f697465723137683765326332623733366531386264656545005f5a4e34636f726533707472376d75745f70747233315f244c5424696d706c2475323024244250246d75742475323024542447542433616464313768333939313037663564323335643062374500497465724d75740047656e657269635261646978006e6578745f696e636c75736976653c636861723e005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243132616c69676e5f6f66667365743137686265366661383332613635626436303545007b696d706c2335337d0064726f705f696e5f706c6163653c26636f72653a3a697465723a3a61646170746572733a3a636f706965643a3a436f706965643c636f72653a3a736c6963653a3a697465723a3a497465723c75383e3e3e005f5a4e34636f7265337074723133726561645f766f6c6174696c653137683034656338646164326362346562306245006d75745f7074720073756d005f5a4e34636f726533666d7439466f726d61747465723770616464696e67313768386664646163386139653836623737364500636d7000696d706c73005f5a4e34636f72653373747232315f244c5424696d706c247532302473747224475424313669735f636861725f626f756e646172793137683034353265303532643135616334353245005f5a4e37355f244c54247573697a65247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c542424753562245424753564242447542424475424336765743137686337356165633633323166633531643545005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542439656e64735f77697468313768383363653331633938643238356662364500696e736572743c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e005f5f72646c5f6f6f6d005f5a4e34636f72653373747235636f756e743131636f756e745f63686172733137683362393037393633646461313835376345007265706c6163653c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e005f5a4e34636f7265366f7074696f6e31354f7074696f6e244c542454244754243769735f736f6d653137686166353061376333383437653666373645006e74683c636f72653a3a7374723a3a697465723a3a43686172496e64696365733e005f5a4e34636f726533737472313176616c69646174696f6e733135757466385f66697273745f627974653137683962396637633933306431356335663945005f5a4e34636f726533666d7438676574636f756e743137683639663830313763343363306364653245005f5a4e34636f72653970616e69636b696e673970616e69635f7374723137683666303932373830653338346562353045005f5a4e34636f726535736c696365366d656d6368723138636f6e7461696e735f7a65726f5f627974653137686130353638656531383330306135373245005f5a4e34355f244c5424244c502424525024247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d74313768613430323766643039663261636331324500666d743c28293e005f5a4e36375f244c5424636f72652e2e61727261792e2e54727946726f6d536c6963654572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d74313768353264643636336235383463633535664500636f70795f6e6f6e6f7665726c617070696e673c75383e00616363756d007b696d706c2334387d007b636c6f7375726523307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542434697465723137686266616536663139613561623764656445006765745f756e636865636b65643c636f72653a3a666d743a3a72743a3a417267756d656e742c207573697a653e006765743c267374723e0070616e69635f646973706c61793c267374723e00756e777261705f6661696c6564002f72757374632f32663662633564323539653761623235646466646433336465353362383932373730323138393138007274005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f7234666f6c64313768623061333862663336373733633236364500636f756e743c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e005f5a4e34636f726533707472347265616431376831653634383335653639376533366630450073756d5f62797465735f696e5f7573697a65005f5a4e34636f726533666d7432727438417267756d656e743861735f7573697a653137686437613231613332353662616362386245005f5a4e3131305f244c5424636f72652e2e697465722e2e61646170746572732e2e656e756d65726174652e2e456e756d6572617465244c54244924475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e657874313768633030313137313163643937383139624500726573756c74005f5a4e37335f244c5424636f72652e2e666d742e2e6e756d2e2e4c6f776572486578247532302461732475323024636f72652e2e666d742e2e6e756d2e2e47656e657269635261646978244754243564696769743137686634306237613733623764393162653445004d61796265556e696e6974007b696d706c2336347d005f5a4e37335f244c54242475356224412475356424247532302461732475323024636f72652e2e736c6963652e2e636d702e2e536c6963655061727469616c4571244c542442244754242447542435657175616c3137686637383434376536346661643333376145005f5a4e3130365f244c5424636f72652e2e6f70732e2e72616e67652e2e52616e6765244c54247573697a6524475424247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c542424753562245424753564242447542424475424336765743137683761383664333261616263343034303345005f5a4e34636f72653463686172376d6574686f647332325f244c5424696d706c247532302463686172244754243131656e636f64655f757466383137683661333732316366346263313738623645005f5a4e34636f726533666d74336e756d33696d7037666d745f7536343137683238366534643532373433386334363745005f5a4e34636f72653970616e69636b696e673570616e69633137686437373538656430613265383739363145006c6962726172792f636f72652f7372632f6c69622e72732f402f636f72652e353431663036343835316338633866372d6367752e3000726561645f766f6c6174696c653c7573697a653e005f5a4e3130385f244c5424636f72652e2e697465722e2e61646170746572732e2e66696c7465722e2e46696c746572244c5424492443245024475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722447542435636f756e7438746f5f7573697a6532385f24753762242475376224636c6f73757265247537642424753764243137686532646263323632336436376436643345005f5a4e34636f726533666d743131506f737450616464696e673577726974653137683130373832303864313037663934393045006164643c7573697a653e005f5a4e34636f726533666d7439466f726d61747465723977726974655f737472313768353330393765363135313339346565644500696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e2c20636f72653a3a6f70733a3a72616e67653a3a52616e676546726f6d3c7573697a653e3e007b696d706c2331357d00656e64735f776974683c75383e005f5a4e34636f726535736c696365366d656d636872366d656d6368723137683838333063653264646237323666636245006c656e5f75746638005f5a4e34636f72653463686172376d6574686f64733135656e636f64655f757466385f7261773137686230336466376165346464366562316445005f5a4e34636f726533666d74355772697465313077726974655f63686172313768666466623438666364333637346132384500616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23347d3a3a6669656c643a3a7b636c6f737572655f656e7623307d3e00636f7265005f5a4e34636f726533636d7035696d706c7335375f244c5424696d706c2475323024636f72652e2e636d702e2e5061727469616c4f72642475323024666f7224753230247573697a6524475424326c74313768383563303932356636663163316566654500646f5f636f756e745f6368617273005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542431336765745f756e636865636b656431376838333832313033623533356331333034450063656c6c006765743c75382c20636f72653a3a6f70733a3a72616e67653a3a52616e67653c7573697a653e3e0066696e6973680077726974655f70726566697800636861725f636f756e745f67656e6572616c5f6361736500706f73745f696e635f73746172743c75383e007265706c6163653c636861723e00506f737450616464696e6700697465723c75383e005f5a4e38375f244c5424636f72652e2e7374722e2e697465722e2e43686172496e6469636573247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683862646365633661316137393933386345005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542433676574313768396431656137353833353464396166364500656e756d6572617465005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683563636236663439653430616432356245005f5a4e34636f726535736c69636534697465723136497465724d7574244c54245424475424336e65773137683131393134666634646337396132326545006469676974005f5a4e34636f726535736c69636533636d7038315f244c5424696d706c2475323024636f72652e2e636d702e2e5061727469616c4571244c54242475356224422475356424244754242475323024666f7224753230242475356224412475356424244754243265713137683331383339323064643563373930336445006d656d6368725f616c69676e656400777261705f6275663c636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23317d3a3a777261703a3a7b636c6f737572655f656e7623307d3e005f5a4e34636f726533666d74386275696c6465727331305061644164617074657234777261703137686630613261643433323636313138356545005f5a4e34636f726533666d74386275696c64657273313044656275675475706c653666696e6973683137683262326465366164386361323965353845006974657200666f6c643c7573697a652c20636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c207573697a652c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e005f5a4e34636f72653373747235636f756e743233636861725f636f756e745f67656e6572616c5f6361736532385f24753762242475376224636c6f73757265247537642424753764243137686238333838383631636166343538396545007b636c6f7375726523307d3c2675382c207573697a652c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e00737065635f6e6578743c7573697a653e005f5a4e34636f726534697465723572616e67653130315f244c5424696d706c2475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722475323024666f722475323024636f72652e2e6f70732e2e72616e67652e2e52616e6765244c5424412447542424475424346e6578743137683166316635393732633862353338396245005f5a4e34636f726533737472313176616c69646174696f6e733138757466385f6163635f636f6e745f62797465313768386431353839303565613233346333334500757466385f6163635f636f6e745f62797465006164643c5b7573697a653b20345d3e006e65773c5b7573697a653b20345d3e005f5a4e34636f726535736c6963653469746572313349746572244c542454244754243134706f73745f696e635f73746172743137686632323465323937613136633263656145006e6578743c636f72653a3a736c6963653a3a697465723a3a497465723c636f72653a3a666d743a3a72743a3a417267756d656e743e3e005f5a4e34636f726535617272617938355f244c5424696d706c2475323024636f72652e2e6f70732e2e696e6465782e2e496e646578244c542449244754242475323024666f722475323024247535622454247533622424753230244e24753564242447542435696e6465783137683663646534633833393961376530333445007b696d706c23397d0064656275675f7475706c655f6e6577005f5a4e34636f726533666d74386275696c64657273313044656275675475706c653666696e69736832385f24753762242475376224636c6f737572652475376424247537642431376861393666623161373161643166373535450064656275675f7475706c655f6669656c64315f66696e697368006164643c75383e007b696d706c233138317d00666f6c643c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a6d61703a3a6d61705f666f6c643a3a7b636c6f737572655f656e7623307d3c2675382c207573697a652c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e3e005f5a4e34636f726535736c69636532395f244c5424696d706c2475323024247535622454247535642424475424313873706c69745f61745f756e636865636b65643137683765396534313435376636393734393145006e6578743c636f72653a3a736c6963653a3a697465723a3a497465723c636f72653a3a666d743a3a72743a3a506c616365686f6c6465723e3e007b696d706c2331377d005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542438697465725f6d75743137683030376635633136366631613761373245006172726179005f5a4e34636f7265337374723469746572323253706c6974496e7465726e616c244c5424502447542431346e6578745f696e636c75736976653137683938613230353930343932666138366445005f5a4e35325f244c542463686172247532302461732475323024636f72652e2e7374722e2e7061747465726e2e2e5061747465726e24475424313269735f7375666669785f6f663137683866653837336364343736333664316445005f5a4e34636f726533666d7439466f726d617474657238777261705f6275663137686636336162363038633262616362303045007b636c6f7375726523307d005f5a4e35365f244c54247573697a65247532302461732475323024636f72652e2e697465722e2e7472616974732e2e616363756d2e2e53756d244754243373756d3137683739356164323965353439386433333445005f5a4e34636f72653373747232315f244c5424696d706c2475323024737472244754243132636861725f696e64696365733137686466343535663065643137623532303045006765743c75382c207573697a653e005f5a4e34636f7265337074723132616c69676e5f6f66667365743137683534623332333739346162326331313545005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243961735f6368756e6b7331376831643562356538303063366463326238450061735f6368756e6b733c7573697a652c20343e005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243361646431376835666664656536393830656665666331450070616e69636b696e67006765745f756e636865636b65643c636f72653a3a666d743a3a72743a3a417267756d656e743e0064656275675f737472756374007b696d706c2332387d0065713c5b75385d2c205b75385d3e0044656275675475706c6500666d745f696e743c636f72653a3a666d743a3a6e756d3a3a55707065724865782c207536343e00636c616e67204c4c564d202872757374632076657273696f6e20312e37312e302d6e696768746c79202832663662633564323520323032332d30352d30392929006974657261746f72005f5a4e34636f726533737472313176616c69646174696f6e7331356e6578745f636f64655f706f696e74313768656364656330303032323838613566354500757466385f66697273745f627974650069735f636861725f626f756e64617279006d696e3c7573697a653e005f5a4e34636f72653373747235636f756e743330636f6e7461696e735f6e6f6e5f636f6e74696e756174696f6e5f627974653137686530636638653465356130663030393045005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137686134633765313364663063343439373145005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243361646431376833356564316564666234363437623138450077726974655f737472005f5a4e34636f726533666d74336e756d313247656e65726963526164697837666d745f696e743137686162643431393537653230363731373445006d617962655f756e696e697400696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e2c20636f72653a3a6f70733a3a72616e67653a3a52616e676546726f6d3c7573697a653e2c203132383e005f5a4e39395f244c5424636f72652e2e7374722e2e697465722e2e53706c6974496e636c7573697665244c54245024475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683536356238663563313134366339666645005f5a4e38315f244c5424636f72652e2e7374722e2e7061747465726e2e2e436861725365617263686572247532302461732475323024636f72652e2e7374722e2e7061747465726e2e2e53656172636865722447542431306e6578745f6d617463683137686231353436643361613035653433333145005f5a4e34636f72653463686172376d6574686f6473386c656e5f75746638313768343935363635353564666635366333654500656e636f64655f757466385f72617700616c6c6f6300747261697473005f5a4e34636f726535736c6963653469746572313349746572244c54245424475424336e65773137683436326338393130346236666239373745005f5a4e34636f7265336e756d32335f244c5424696d706c24753230247573697a652447542431327772617070696e675f6d756c3137683933396664623563663661656266303945006e6577006d656d6368720077726170005f5a4e34636f726533666d74336e756d313247656e65726963526164697837666d745f696e743137683330323730653937613764383866626145007061640070616e6963005f5a4e34636f726533666d74336e756d35335f244c5424696d706c2475323024636f72652e2e666d742e2e4c6f7765724865782475323024666f7224753230246936342447542433666d74313768663235653065383534373535336437314500696d7000616c7465726e617465006d6170005f5a4e3130325f244c5424636f72652e2e697465722e2e61646170746572732e2e6d61702e2e4d6170244c5424492443244624475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722447542434666f6c643137683439653563633739303661396231626645007772697465007b696d706c23377d006d696e5f62793c7573697a652c20666e28267573697a652c20267573697a6529202d3e20636f72653a3a636d703a3a4f72646572696e673e006765743c267374722c207573697a653e005f5a4e34636f726535736c69636535696e64657837345f244c5424696d706c2475323024636f72652e2e6f70732e2e696e6465782e2e496e646578244c542449244754242475323024666f72247532302424753562245424753564242447542435696e64657831376835623336343435386238326632343635450053706c6974496e7465726e616c006e6578743c636861723e0057726974650077726974655f636861723c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e007b696d706c2332367d005f5a4e34636f72653970616e69636b696e67313870616e69635f6e6f756e77696e645f666d743137683133386130386530383963323036303445005f5a4e34325f244c54242452462454247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d74313768633230363132656137383639386165344500666d74007b696d706c23307d004f7074696f6e007b696d706c23387d005f5a4e34636f726533707472376d75745f70747233315f244c5424696d706c2475323024244250246d757424753230245424475424336164643137686433383935323761353331303836366545006765745f756e636865636b65643c267374723e005f5a4e34636f726533666d7439466f726d6174746572313264656275675f73747275637431376838333134343030643138313466376534450070616e69635f737472005f5a4e34636f726533666d74386275696c64657273313564656275675f7475706c655f6e65773137683134383664383033383865636636373745005553495a455f4d41524b455200736c696365005f5a4e34636f7265336d656d377265706c6163653137683665313530623565366261663964346545007061645f696e74656772616c006765743c75383e005f5a4e34636f726535736c6963653469746572313349746572244c54245424475424336e65773137686231373834333338323430613463363745007b696d706c2331397d006e6578745f6d61746368005f5a4e34636f726536726573756c743139526573756c74244c542454244324452447542438616e645f7468656e3137686639613762303833656534636237383245005f5a4e37335f244c5424636f72652e2e666d742e2e6e756d2e2e5570706572486578247532302461732475323024636f72652e2e666d742e2e6e756d2e2e47656e657269635261646978244754243564696769743137683933663339316566393536306361643245005f5a4e34636f72653370747231303264726f705f696e5f706c616365244c542424524624636f72652e2e697465722e2e61646170746572732e2e636f706965642e2e436f70696564244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c542475382447542424475424244754243137683465633534623435323134663763393045005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683334323336653433336537396333623345006c74006368617273005f5a4e34636f72653373747232315f244c5424696d706c247532302473747224475424336765743137686361316261643162613538333362626645006765743c636f72653a3a6f70733a3a72616e67653a3a52616e6765546f3c7573697a653e3e00706f73745f696e635f73746172743c7573697a653e005f5a4e37355f244c54247573697a65247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c54242475356224542475356424244754242447542431336765745f756e636865636b65643137686630663432666234656339376261626145006164643c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e006d6574686f6473005f5a4e34636f726533666d74386275696c64657273313050616441646170746572347772617032385f24753762242475376224636c6f737572652475376424247537642431376862353032353031383864353564626337450063617061636974795f6f766572666c6f7700666d745f753634005f5a4e36385f244c5424636f72652e2e666d742e2e6275696c646572732e2e50616441646170746572247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f7374723137686539366438303337316562386433343445005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243361646431376836343831303738333031643161616237450049746572005f5a4e34636f72653373747232315f244c5424696d706c2475323024737472244754243563686172733137683635643537336338666664393434333645005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f723130616476616e63655f62793137683837343136383366376333383664636245006e6578745f636f64655f706f696e743c636f72653a3a736c6963653a3a697465723a3a497465723c75383e3e005f5a4e39335f244c5424636f72652e2e736c6963652e2e697465722e2e4368756e6b73244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137686264343939663734373230663065386245004f7264006164643c267374723e007b696d706c23367d005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f666d743137683565373464633863623261616161323645007b696d706c23327d005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542434697465723137686331616261316236653465646465623545005f5a4e34636f726533666d7439466f726d6174746572336e65773137686165623034366666366431666231663445005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243361646431376838353436653232346135313966363633450064656275675f7374727563745f6e657700746f5f7538005f5a4e34636f726533636d7035696d706c7336395f244c5424696d706c2475323024636f72652e2e636d702e2e5061727469616c4571244c54242452462442244754242475323024666f7224753230242452462441244754243265713137683436393566636435376362636161326145005f5a4e34636f726533666d743577726974653137683537653362636463656237646630393145006578706563745f6661696c6564006c656e5f6d69736d617463685f6661696c006f707300696e7472696e736963730073756d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e005f5a4e34636f7265336d656d377265706c61636531376838363534306363336630326138396663450069735f6e6f6e653c7573697a653e00697465723c5b7573697a653b20345d3e00696e746f5f697465723c5b7573697a653b20345d3e005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683366313636623661373436326234373945005f5a4e34636f726533666d7432727438417267756d656e7433666d74313768363232636537653835383430326338654500666d745f696e743c636f72653a3a666d743a3a6e756d3a3a4c6f7765724865782c207536343e00657175616c3c75382c2075383e005f5a4e34636f726535736c696365366d656d63687231326d656d6368725f6e616976653137686363623962373463393862393633336245006d656d6368725f6e6169766500616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23347d3a3a66696e6973683a3a7b636c6f737572655f656e7623307d3e005f5f616c6c6f635f6572726f725f68616e646c657200636f6e73745f707472005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f723373756d313768616537613566613764646461346162384500757466385f69735f636f6e745f62797465006e6578743c636f72653a3a666d743a3a72743a3a417267756d656e743e005f5a4e34636f726533666d74386275696c64657273313664656275675f7374727563745f6e65773137686135363836656238343531653037323245005f5a4e34636f72653970616e69636b696e67313370616e69635f646973706c6179313768663965353336303933393038663832624500656e64735f776974683c636861723e0065713c75382c2075383e007b696d706c23347d005f5a4e34636f726533737472313176616c69646174696f6e733137757466385f69735f636f6e745f6279746531376861396331376363326537313134623836450073706c69745f61745f756e636865636b65643c75383e0073706c69745f61743c75383e005f5a4e34636f72653373747235636f756e74313873756d5f62797465735f696e5f7573697a653137683733663965326535343130353136333245006e6578743c636f72653a3a666d743a3a72743a3a506c616365686f6c6465723e00417267756d656e74005f5a4e37355f244c54247573697a65247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c54242475356224542475356424244754242447542431336765745f756e636865636b6564313768656630633435353430343632353962624500636f6e7461696e735f7a65726f5f62797465005f5a4e37395f244c5424636f72652e2e726573756c742e2e526573756c74244c5424542443244524475424247532302461732475323024636f72652e2e6f70732e2e7472795f74726169742e2e54727924475424366272616e63683137683034646133323232663535363066313845005f5a4e34636f7265366f7074696f6e31336578706563745f6661696c65643137686332333330616533386638616564396545005f5a4e34636f726533707472376d75745f70747233315f244c5424696d706c2475323024244250246d7574247532302454244754243361646431376837336363316163653933303039363536450073756d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e2c207573697a653e005f5a4e35365f244c54247573697a65247532302461732475323024636f72652e2e697465722e2e7472616974732e2e616363756d2e2e53756d244754243373756d32385f24753762242475376224636c6f73757265247537642424753764243137683665653564323561643365666465373945007369676e5f61776172655f7a65726f5f70616400726561643c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e006e6578743c7573697a653e00756e777261705f6f723c267374723e005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243136616c69676e5f746f5f6f6666736574733137683265333033653231353164623038353745005f5a4e34636f726535736c69636532395f244c5424696d706c2475323024247535622454247535642424475424336765743137683037666466393631613031323632356145006e65773c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e007b696d706c2334347d0070616e69635f6e6f756e77696e645f666d740077726974655f7374723c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e577269746524475424313077726974655f636861723137683239666437616639333939643762333645005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243135636f70795f66726f6d5f736c69636531376c656e5f6d69736d617463685f6661696c3137686531663934356265353831313135613845006c6962726172792f616c6c6f632f7372632f6c69622e72732f402f616c6c6f632e643733613839653266303538366464312d6367752e30004974657261746f7200636f756e745f6368617273005f5a4e34636f72653469746572386164617074657273336d6170386d61705f666f6c6432385f24753762242475376224636c6f73757265247537642424753764243137686265643362346664336632356561633645005f5a4e34636f7265366f7074696f6e31354f7074696f6e244c542454244754243769735f6e6f6e653137683036303537623832613939663564313445005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542438616c69676e5f746f3137686361663565313535373365303734303345007b696d706c2331317d005f5a4e34636f726533636d70366d696e5f62793137683961363365346463336265666132393045005f5a4e34636f7265336d656d31326d617962655f756e696e697432304d61796265556e696e6974244c54245424475424357772697465313768643262633963366561386361383161624500656e636f64655f75746638005f5a4e34636f726533666d743557726974653977726974655f666d743137683364623431343565346436363932376245006669656c64005f5a4e36305f244c5424636f72652e2e63656c6c2e2e426f72726f774572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137686163386261333334363731373261333845006e6578743c75383e00746f5f7573697a65006d656d005f5a4e34636f7265337074723577726974653137683934303032343231393363646338316545005f5a4e38395f244c5424636f72652e2e6f70732e2e72616e67652e2e52616e6765244c54245424475424247532302461732475323024636f72652e2e697465722e2e72616e67652e2e52616e67654974657261746f72496d706c2447542439737065635f6e65787431376834303038636235396134653064623339450061735f7573697a65006164643c636f72653a3a666d743a3a72743a3a417267756d656e743e00696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e005f5a4e34636f7265336e756d32335f244c5424696d706c24753230247573697a652447542431327772617070696e675f73756231376838643635306338643866353735643162450069735f70726574747900616461707465727300726561643c636861723e007b696d706c23337d00636861725f696e646963657300616c69676e5f746f3c75382c207573697a653e007772617070696e675f6d756c0077726974653c75383e005f5a4e35305f244c5424753634247532302461732475323024636f72652e2e666d742e2e6e756d2e2e446973706c6179496e742447542435746f5f75383137683636316463333963356464386666653545007061747465726e0069735f7375666669785f6f66005f5a4e34636f726535736c696365366d656d63687231346d656d6368725f616c69676e6564313768643864383232303663636532343531614500526573756c740050616441646170746572005f5a4e34636f726533666d7439466f726d6174746572337061643137683433336537613934646232626438653245005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f7374723137683865303931326361326264646233386345005f5a4e34636f726533666d7432727431325553495a455f4d41524b455232385f24753762242475376224636c6f7375726524753764242475376424313768643137376134333532613130653633314500466e4f6e6365006e756d005f5a4e38315f244c5424636f72652e2e7374722e2e697465722e2e4368617273247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722447542435636f756e743137686638633866336432633063356164333545005f5a4e34636f726533666d7439466f726d617474657231397369676e5f61776172655f7a65726f5f7061643137683136323439616566366630343733333545006e65773c75383e007b696d706c23357d005f5a4e34636f726533636d70334f7264336d696e31376861623865636338303366663033636364450072756e005f5a4e34636f726533666d74386275696c64657273313044656275675475706c653969735f7072657474793137683131646663373739346165376162303045005f5a4e34636f726533666d7439466f726d617474657231327061645f696e74656772616c313277726974655f70726566697831376838346635386564303837613362643933450066756e6374696f6e00466f726d61747465720066696c746572006d61705f666f6c64005f5a4e38315f244c5424636f72652e2e7374722e2e697465722e2e4368617273247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683064323235303663643135633337363345007b696d706c2337307d005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683634663237353939353136663335636545005f5a4e35355f244c542424524624737472247532302461732475323024636f72652e2e7374722e2e7061747465726e2e2e5061747465726e24475424313269735f7375666669785f6f663137686536396533336230613062663235373545007772617070696e675f7375620077726974655f666d743c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e005f5a4e35616c6c6f63377261775f766563313763617061636974795f6f766572666c6f7731376837363964333737343539393364316265450063616c6c5f6f6e63653c636f72653a3a666d743a3a72743a3a5553495a455f4d41524b45523a3a7b636c6f737572655f656e7623307d2c2028267573697a652c20266d757420636f72653a3a666d743a3a466f726d6174746572293e0062000000020000000000740000003400000063617061636974795f6f766572666c6f77002f0000007261775f76656300590000005f5f72646c5f6f6f6d004f000000616c6c6f6300540000005f5f616c6c6f635f6572726f725f68616e646c65720000000000de1a0000020074000000cb2200006a01000077726974653c636861723e00c61e00006d617962655f756e696e6974007c2100006272616e63683c28292c20636f72653a3a666d743a3a4572726f723e00e90000006d75745f707472008a1f0000696e736572743c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e0003190000636f70795f6e6f6e6f7665726c617070696e673c75383e00b7040000466f726d617474657200752000007b696d706c2331377d00b01c0000737065635f6e6578743c7573697a653e0086190000706f73745f696e635f73746172743c7573697a653e00381800007b696d706c2332357d0057210000526573756c7400cb1d00006e6578745f636f64655f706f696e743c636f72653a3a736c6963653a3a697465723a3a497465723c75383e3e0034000000726561645f766f6c6174696c653c7573697a653e002b1a0000697465723c5b7573697a653b20345d3e00b91e00007265706c6163653c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e00711c00007b636c6f7375726523307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e00f719000073706c69745f61745f756e636865636b65643c75383e00ac1e00007265706c6163653c636861723e00701f000069735f6e6f6e653c7573697a653e00451a00006765743c267374722c207573697a653e00b02100007b696d706c2332367d00271e000069735f636861725f626f756e646172790038210000726573756c74008718000066756e6374696f6e00671c0000636f756e7400f00400007061645f696e74656772616c00111a0000616c69676e5f746f5f6f6666736574733c75382c207573697a653e008b1a00006c656e5f6d69736d617463685f6661696c00da0000006164643c75383e006e1900006e65773c75383e00e203000064696769740050180000666d743c28293e001f20000070616e69636b696e67007d1f0000756e777261705f6f723c267374723e00451d0000636f6e7461696e735f6e6f6e5f636f6e74696e756174696f6e5f6279746500cd000000616c69676e5f6f66667365743c75383e00bd1900006e65773c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e00d62000007b696d706c2331397d00102000007772617070696e675f73756200c9040000616c7465726e61746500fc1e00006c74003e1c00006d61705f666f6c6400511d000073756d5f62797465735f696e5f7573697a6500ae010000417267756d656e7400cb1e00004d61796265556e696e697400f4030000666d7400981f00006578706563745f6661696c6564009f1b0000636f6e7461696e735f7a65726f5f6279746500a911000072756e00a61d00007b696d706c2334347d006c1e00007b696d706c2332387d008d11000077726974655f707265666978008c180000466e4f6e636500d61a00006765743c267374723e005b000000636f6e73745f70747200971e00006e6578745f6d6174636800791a00006765743c75382c20636f72653a3a6f70733a3a72616e67653a3a52616e67653c7573697a653e3e00dd1e000077726974653c75383e00340100006164643c7573697a653e005d19000049746572003713000064656275675f7374727563745f6e6577004b1800007b696d706c2335337d00b30000006164643c636f72653a3a666d743a3a72743a3a417267756d656e743e00ed1c0000737472003d20000070616e69635f646973706c61793c267374723e00d0190000697465723c75383e00861a0000636f70795f66726f6d5f736c69636500271c00006d617000671e00007061747465726e00d9020000666d745f696e743c636f72653a3a666d743a3a6e756d3a3a4c6f7765724865782c207536343e00b015000066696e69736800dd0300007b696d706c2332397d0069210000616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23347d3a3a66696e6973683a3a7b636c6f737572655f656e7623307d3e003d210000756e777261705f6661696c656400201900006e6578743c75383e00931d000053706c6974496e7465726e616c00211d0000646f5f636f756e745f636861727300501900006e6578743c636f72653a3a666d743a3a72743a3a417267756d656e743e0011190000736c69636500c415000044656275675475706c65006c1c0000746f5f7573697a650062190000706f73745f696e635f73746172743c75383e005e1d000069746572000d1c000073756d00f71e00007b696d706c2335347d00931900007b696d706c2337307d00ca1a00006765745f756e636865636b65643c636f72653a3a666d743a3a72743a3a417267756d656e743e00841700007b696d706c23307d000f1d0000636861725f636f756e745f67656e6572616c5f6361736500841e000069735f7375666669785f6f6600311c0000666f6c643c7573697a652c20636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c207573697a652c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e007f100000777261705f6275663c636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23317d3a3a777261703a3a7b636c6f737572655f656e7623307d3e000918000077726974655f666d743c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e00e3010000666d745f753634002a000000636f7265001e1a000061735f6368756e6b733c7573697a652c20343e006211000064656275675f7475706c655f6669656c64315f66696e697368009c0100005553495a455f4d41524b455200221c0000616461707465727300f61f00007772617070696e675f6d756c00121c00007b636c6f7375726523307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e00331e00006765743c636f72653a3a6f70733a3a72616e67653a3a52616e6765546f3c7573697a653e3e00a60000006164643c5b7573697a653b20345d3e005b1c0000636f756e743c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e00ab190000696e746f5f697465723c5b7573697a653b20345d3e00c11b0000666f6c643c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a6d61703a3a6d61705f666f6c643a3a7b636c6f737572655f656e7623307d3c2675382c207573697a652c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e3e00e11600007b696d706c23317d005520000070616e69635f6e6f756e77696e645f666d7400902200006368617200511c000066696c74657200811c0000656e756d6572617465007b1b00006d656d6368725f6e6169766500e304000070616464696e6700160300007b696d706c2336347d00fc1b00007b696d706c2334387d00e61600007772617000f916000064656275675f7475706c655f6e657700431300007b696d706c23327d00b301000061735f7573697a6500011c000073756d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e00f21e0000696d706c7300f71b0000616363756d00071700005772697465002420000070616e696300441900006e6578743c636f72653a3a666d743a3a72743a3a506c616365686f6c6465723e000d1e0000636861727300821800006f707300952200006d6574686f6473005c1b000065713c75382c2075383e00ab1d00006e6578743c636861723e00ef0300007b696d706c2336357d00401e0000656e64735f776974683c636861723e00a71e00006d656d007f1e00007b696d706c23337d004920000070616e69635f73747200d61500006669656c6400381f00004f72640097010000727400de010000696d70008b1c00006e6578743c636f72653a3a736c6963653a3a697465723a3a497465723c636f72653a3a666d743a3a72743a3a506c616365686f6c6465723e3e00381900006e6578743c7573697a653e00b8190000497465724d757400c31100007772697465005f1a0000656e64735f776974683c75383e00c915000069735f707265747479002c1900006e6578743c5b7573697a653b20345d3e00e5020000666d745f696e743c636f72653a3a666d743a3a6e756d3a3a55707065724865782c207536343e00db1b0000616476616e63655f62793c636f72653a3a7374723a3a697465723a3a43686172496e64696365733e00d402000047656e657269635261646978004e1e0000747261697473008917000077726974655f7374723c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e00861d00006e65787400ce1b000073756d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e2c207573697a653e00981500007b696d706c23347d004813000077726974655f737472009a2200006c656e5f75746638001c1f000065713c5b75385d2c205b75385d3e005d010000726561643c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e00041a000073706c69745f61743c75383e00981d00006e6578745f696e636c75736976653c636861723e00040300007b696d706c2331317d0050010000726561643c636861723e00d907000070616400431c00007b636c6f7375726523307d3c2675382c207573697a652c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e00a217000077726974655f636861723c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e00d71d0000757466385f66697273745f6279746500391b00007b696d706c23357d00971c00006e6578743c636f72653a3a736c6963653a3a697465723a3a497465723c636f72653a3a666d743a3a72743a3a417267756d656e743e3e002b1f00006d696e5f62793c7573697a652c20666e28267573697a652c20267573697a6529202d3e20636f72653a3a636d703a3a4f72646572696e673e00591000006e657700df1f00006e756d007701000077726974653c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e00b41a0000696e646578005e1f00004f7074696f6e00631f000069735f736f6d653c7573697a653e00321300006275696c64657273001a1e0000636861725f696e6469636573007020000063656c6c00c00000006164643c267374723e00dd1900006765743c75382c207573697a653e00ef1a00007b696d706c23367d00251b00006765743c75383e00b51500007b636c6f7375726523307d00bf1d0000757466385f69735f636f6e745f6279746500bc1b00004974657261746f72009118000063616c6c5f6f6e63653c636f72653a3a666d743a3a72743a3a5553495a455f4d41524b45523a3a7b636c6f737572655f656e7623307d2c2028267573697a652c20266d757420636f72653a3a666d743a3a466f726d6174746572293e00871b00006d656d6368725f616c69676e656400ea190000616c69676e5f746f3c75382c207573697a653e00381a00006765745f756e636865636b65643c636f72653a3a666d743a3a72743a3a417267756d656e742c207573697a653e00410100006164643c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e00a61a0000697465725f6d75743c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e00591f00006f7074696f6e00a7220000656e636f64655f757466385f72617700ba1d000076616c69646174696f6e7300341b0000636d7000581e000067657400e21a00006765745f756e636865636b65643c267374723e00831100007b696d706c23377d001b1900007b696d706c233138317d00b71b00006974657261746f72007210000064656275675f73747275637400131b0000696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e2c20636f72653a3a6f70733a3a72616e67653a3a52616e676546726f6d3c7573697a653e3e00e81b00006e74683c636f72653a3a7374723a3a697465723a3a43686172496e64696365733e00b9220000656e636f64655f7574663800cf16000050616441646170746572006f1b00006d656d63687200531e00007b696d706c23387d00d7180000696e7472696e7369637300a2210000696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e2c20636f72653a3a6f70733a3a72616e67653a3a52616e676546726f6d3c7573697a653e2c203132383e00a61c000072616e676500902100007b696d706c2331357d00d60400007369676e5f61776172655f7a65726f5f70616400bc0400007369676e5f706c7573002f000000707472004100000064726f705f696e5f706c6163653c26636f72653a3a697465723a3a61646170746572733a3a636f706965643a3a436f706965643c636f72653a3a736c6963653a3a697465723a3a497465723c75383e3e3e00031d0000636f756e745f6368617273007a1900006e65773c5b7573697a653b20345d3e0070110000506f737450616464696e6700fb1d0000757466385f6163635f636f6e745f6279746500f41a0000696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e000a1f00007b696d706c23397d00b6110000676574636f756e74005c210000616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23347d3a3a6669656c643a3a7b636c6f737572655f656e7623307d3e004b1f00006d696e3c7573697a653e0009030000746f5f7538003e1b0000657175616c3c75382c2075383e008b210000617272617900000000000e00000002000000000074000000000000000e000000020074000000cb22000000000000412a000000726973637600012000000004100572763634693270305f6d3270305f613270305f633270300084000000040040000000010101fb0e0d0001010101000000010000016c6962726172792f616c6c6f632f73726300007261775f7665632e727300010000616c6c6f632e727300010000000009029a42010000000000038a040105050a030109020001090c000001010402000902a842010000000000038d0301050d0a030b09020001090c00000101ed1b0000040052030000010101fb0e0d0001010101000000010000016c6962726172792f636f72652f7372632f6f7073006c6962726172792f636f72652f7372632f707472006c6962726172792f636f72652f7372632f666d74006c6962726172792f636f72652f737263006c6962726172792f636f72652f7372632f736c6963652f69746572006c6962726172792f636f72652f7372632f697465722f747261697473006c6962726172792f636f72652f7372632f737472006c6962726172792f636f72652f7372632f69746572006c6962726172792f636f72652f7372632f697465722f6164617074657273006c6962726172792f636f72652f7372632f6d656d006c6962726172792f636f72652f7372632f6d6163726f73006c6962726172792f636f72652f7372632f736c696365006c6962726172792f636f72652f7372632f6e756d006c6962726172792f636f72652f7372632f6172726179006c6962726172792f636f72652f7372632f63686172000066756e6374696f6e2e7273000100006d6f642e72730002000072742e7273000300006e756d2e727300030000636f6e73745f7074722e727300020000696e7472696e736963732e7273000400006d75745f7074722e7273000200006d6f642e7273000300006d6163726f732e7273000500006974657261746f722e72730006000076616c69646174696f6e732e727300070000616363756d2e727300060000636d702e72730004000072616e67652e7273000800006d61702e72730009000066696c7465722e727300090000636f756e742e727300070000697465722e7273000700006d6f642e7273000a00006f7074696f6e2e7273000400006d6f642e7273000b00006d6f642e727300070000696e6465782e7273000c00007472616974732e7273000700006d6f642e7273000c000075696e745f6d6163726f732e7273000d0000697465722e7273000c000070616e69636b696e672e727300040000656e756d65726174652e72730009000063656c6c2e7273000400006275696c646572732e727300030000726573756c742e7273000400006d617962655f756e696e69742e7273000a00006d6f642e7273000e0000636d702e7273000c00007061747465726e2e7273000700006d656d6368722e7273000c00006d6574686f64732e7273000f000000000902747701000000000003f90101040205090a03860a090000010403050503d375090200010902000001010402000902787701000000000003ea030105010a03000900000109020000010104040009027a7701000000000003d2010105170a03130906000106039a7e0918000103e60109040001039a7e0924000105150603e80109020001051e0302090e00010405050d03b505091a00010406050903d20d090200010404051e03fa6c0904000104060509038613090400010405050d03ae72090800010406050903d20d090200010404051503fb6c09080001040605090385130902000106030009040001040405170603f56c0908000106039a7e0906000105140603f901090400010515030209040001051e037f091c000105150302090400010405050d03a305090200010406050903d20d090200010407050d039c73090c00010406050903e40c0902000106038f6b090a000104040514060381020902000105150301090400010407050d038b06090800010404051503f67909020001051e0302090a000105150301090200010405050d039905090400010406050903d20d090200010407050d039c73090c00010406050903e40c0902000106038f6b090800010407050d06038d08090400010404053e03827a09060001050d030209020001050a030109140001060b0300090200010904000001010408000902bc7801000000000003dd090105090a03e003091e0001051303a77c090c000106039b76090c000105090603f70d09040001051303ee7b0904000105190305090200010603967609020001050f0603fb0909020001050906030009020001038576090400010409051806038601090200010603fa7e09040001040a05150603b113090400010407050d03dc7409040001040b0505038c78090200010409051803ed0009080001040c051c03af7f090200010409051803d100090200010408050d03e50809020001050f031009020001050906030009020001052306030909020001051a06030009040001050906038d0409040001051a03f97b09020001051b03e90009020001053103a47f09060001051503dc000904000106038d7509060001050606039d0a09200001060b0300091c0001050003e3750904000104020509060394090926000106030009060001040805110603f900090400010402050903cd00090a000106030009040001040805110603b37f090400010603f3750914000105090603800b09020001040d05340353090600010408050d032e090400010603ff740910000105150603f30a090200010530030a0904000105230603000904000105300300090200010383750906000105090603800b090c0001040d0534035309040001040e050c039a7a090200010408050d039406090200010603ff74090c000105240603970a090a00010511030109040001030109140001050903fb7e090e0001040d053403bf01090800010408050d03c27e09080001051103fa00091000010603f175091000010603910a090200010301090400010603ee7509080001040d05340603d30a090200010906000001010408000902a07a01000000000003f2090105140a0301091c0001051103010904000105140302090e0001052c060300090200010b03000912000103897609040001050a0603f80909020001060b0300090a00010904000001010408000902f67a01000000000003bb0a01041405120a039b7a090200010408050c03e7050916000104150509039a78090200010408050c03e607090800010518030509040001051d060300090400010405050d0603dc7c09040001040a050903b87b09040001040b05000603a97d09120001041205260603910109040001051106030009020001040a05100603c70109040001040d053403fb0709040001040e050c039a7a090200010409051803997c09020001040b050d03a07f0904000105080301090800010516030a090400010505035b0904000105110306090400010508032109040001051a0305090400010505035a090400010511060300090200010505030009040001050c06032909040001051e030509040001051203010904000105050351090400010511060300090200010505030009040001050d06032f090400010412050903cb00090200010603f47e090400010409051806038601091e0001040b050d03a07f090400010508030109040001060359090400010603330908000106034d09040001050c06033b09040001050006034509040001051a060338090400010511035a0904000106030009040001051e06032e09040001051203010904000105050351090400010511060300090600010505030009040001050d06032f090200010412050903cb00090600010416050c03cc000904000105090304090200010417050c037d0904000104160513030f0904000104180509032c090800010603ec7d0904000104140603bc0709020001041803d87a090400010603ec7d0904000104140603bc07090200010603c4780902000104080603d40a0904000105120304090400010411050803c37509080001060365090400010409051806038601090200010603fa7e09040001040a05150603b113090400010407050d03dc7409040001040b0505038c78090200010409051803ed0009080001040c051c03af7f090200010409051803d100090200010402051f03bb0c0904000104190545036509060001051603800e090800010409051803e065090600010603fa7e09040001040a05150603b113090200010407050d03dc7409040001040b0505038c78090200010409051803ed0009080001040c051c03af7f090200010409051803d100090200010603fa7e090200010386010902000103fa7e09020001040a05150603b113090600010407050d03dc7409040001040b0505038c78090200010409051803ed0009080001040c051c03af7f090200010409051803d100090200010603fa7e09020001041105150603c7000922000105000603b97f09060001051b0603fe00090e00010534060300090400010533030009020001051b030009040001041a050d0603e7080902000104110505039a77090400010509035b09020001050c030609020001041b03e80a090200010603b874090200010419053806039908091200010405050d03867f090400010409051803e779090600010603fa7e09020001041105190603d0000904000105120301090200010507032309020001050606030009040001051203000902000106035d09020001050503230902000105110360090400010507032009020001050606030009040001051206035d090200010323090200010505060300090200010507030009040001050603000904000105120300090200010505030009020001051206035d0902000105050323090200010511036009020001050703200904000105060603000904000105120300090200010505030009020001040905180603120904000104110511034e09040001040905180332090200010603000906000103fa7e090400010386010904000103fa7e09040001038601090600010411051206035d090600010407050d03aa07090200010411050703e7780902000105060603000904000105120300090200010505030009020001040905180603120904000104110511035e09020001040905180322090200010603fa7e090400010411051b0603fe00090200010534060300090400010533030009020001051b030009040001041a050d0603e7080902000104110505039a7709040001050d0367090200010408051403f60909020001051b0317090400010535037009060001051503100904000106038d750906000103f30a09260001053006030a0904000105230603000904000105300300090200010383750906000105090603800b090e0001040d0534035309040001040e050c039a7a090200010408050d039406090200010603ff74090c000105280603e30a090a00010515030109040001050903b07e090e0001040d053403bf0109080001040e050c039a7a090400010408050d03a804090400010603eb7609100001040d05340603d30a0902000104080506031609040001060b030009140001090400000101041c0009026e7e01000000000003ed000105050a030709020001090c0000010104080009027c7e01000000000003b7080105090a03bb7909180001050b03c90609080001050903b77909040001050503c90609080001050e030e090200010409051803bc78090400010603fa7e0904000103860109040001040805150603cb0709220001051406030009020001051506030109020001052d0603000904000105150300090400010510060313090600010505060300090200010511060301090200010505060300090400010511060301090400010533036f09020001050503110904000105150304090200010505030f090600010403050c039978090600010603ed7e090a0001051d0603960109040001051b0603000902000103ea7e09020001040805090603eb080902000105190301090400010505030e090800010403050c039978090600010603ed7e090a0001051d0603960109040001051b0603000902000103ea7e09020001040805090603ec0809020001052d0307090400010405050d03ac7e090200010403050903eb7909040001051a060300090200010509030009020001040805110603cc07090400010409051803b078090200010408051d03b907091000010409051803c778090400010603fa7e0904000103860109080001040805150603bd0709120001051406030009020001051506030109020001052d060300090400010515030009040001040305090603c67809060001051a060300090200010509030009040001040805110603bc07090400010409051803c078090200010408051a03d707090a00010417050c03fc78090400010603a77e090600010408051a0603dd08090200010417050c03fc78090400010408051a038407090400010405050d03c27e090400010408050903bf0109040001052106030009040001050903000908000103a2770906000105020603e20809060001060b030009100001090400000101041e000902fa7f01000000000003ba0501040805090a03ba0609000001091200000101041e0009020c8001000000000003d50501040805090a039f060900000109120000010104200009021e8001000000000003f10c0105050a030109020001090c0000010104140009022c80010000000000038a0f01041c05050a038b7209020001090c00000101041c0009023a8001000000000003cf0001050e0a031009020001090c0000010104040009024880010000000000039901010407050d0a03f30609060001040405000603f3770908000106039301090800010421050903d602090200010404051403ea7c090400010603ad7f09080001052306032a0902000103e900090800010603ed7e090400010417050c0603ed03090a00010404050903817d090a0001050e032e09160001060b0300090200010417050d0603d20209040001090e00000101041f000902b880010000000000031e010412050c0a03ce040946000104190523039c0d091800010423050d03d26e09040001041f034a090a00010301090400010412050c03c704090e00010424051903b17e090800010417050c0342090a00010425050803cb7d09080001050b030d0906000106034809040001050c0603390902000105090304090c0001050b037b090200010402051f03890d09060001051b03010908000104250508039273090400010603ac7f090e000105100603eb00090600010405050d03b406090400010425051503c679090400010529030409060001041a050d03e508090200010425050503c67609020001051503d2000908000105290304090a0001041a050d03e408090200010425050503c67609020001050903db0009080001050b037209020001050c03580906000105090304090c0001050b037b09020001060348090400010603e1000904000106039f7f09040001050c06033909060001050b037f090c000106034809080001042405200603b403090200010511060300090200010417050c0603ac7f090800010423050d03fb7d090200010424051c03dd02090400010603c87c09040001041f051006032109140001051103010906000106035e090e00010419050906038912090800010603f76d09040001041f050606032a09100001060b0300091a00010904000001010408000902748201000000000003a20101052b0a0301090c00010426050803f60b09020001050d031f09040001050f0363090800010513032009060001050d06030009040001051206030109080001050d06030009040001050f060361090c00010513032209060001050d06030009040001051206030109080001050d06030009060001051206030109080001050d060300090400010512060303090c0001050d06030009060001051206030109080001050d06030009060001051206030109080001050d06030009060001051206030109080001050d06030009040001040805090603dc73090a000105060301090a0001060b0300090200010904000001010408000902288301000000000003be010105090a0301090200010506030109300001060b0300090200010904000001010408000902608301000000000003c5010105090a030109000001090a0000010104080009026a8301000000000003c9010105090a030109020001052b0359090c00010426050803f60b09020001050d031f09040001050f0363090800010513032009060001050d06030009040001051206030109080001050d06030009040001050f060361090c00010513032209060001050d06030009040001051206030109080001050d06030009060001051206030109080001050d060300090400010512060303090c0001050d06030009060001051206030109080001050d06030009060001051206030109080001050d06030009060001051206030109080001050d06030009040001040805090603dc73090a000105060328090a0001060b0300090200010904000001010408000902208401000000000003cd010105090a0301090200010371091e00010506031009140001060b030009020001090400000101041f0009025a8401000000000003b3020105170a0301091200010420050903f10709040001041f03a078090200010603ba7d0908000105100603b602090400010408050903c10b09040001041f050006038972090400010408050903f70d09040001041f05100603bf740904000105000603ca7d09020001051e0603c002090400010603c07d0904000105140603b702090a00010408050903be0909040001041f051503c376091600010603c87d09020001040805090603f50b090e0001041f051e03cb76090a00010408050903b50909020001042003a70309040001041f051103a673090200010408051403e406090c00010603da7609040001041f05210603bb02090200010408051703e806090400010414050903f002090800010408051303947d090a0001051403010904000103010904000105180301090800010509037709080001041f0511039c79091400010408050903e40609040001041f0511039c79090a00010408050903b80909080001041f050006038b740912000105090603b502090200010311090400010506030209060001060b03000910000109040000010104080009027a8501000000000003e40f0105090a03907c090c0001041f050503a376090c00010408050903cf0d090c0001041f050c03fd72090e0001050006039c7d09020001050c03e40209040001039c7d09020001042005090603a60a09020001041f051403c07809020001050006039a7d090a0001051403e60209020001040805090603910b09080001041f051403ef740906000104080509038f0909020001041f051503f2760914000104080509038e0909020001041f03f776091600010408050603fd0c09040001060b0300090a000109040000010104190009021286010000000000038a1a01050d0a030109020001090c000001010408000902208601000000000003cf110105090a03ec01090000010916000001010422000902368601000000000003820101040805090a03f20a090a00010422051e038f75090200010408050903f10a09020001041f050503a376091000010408050903cf0d090c0001041f050c03fd7209140001050006039c7d09020001050c03e40209040001039c7d09020001042005090603a60a09020001041f051403c07809020001050006039a7d090a0001051403e60209020001040805090603910b09080001041f051403ef740906000104080509038f0909020001041f051503f2760914000104080509038e0909020001041f03f776091600010422050f03977e09040001060b0300090800010904000001010404000902d886010000000000039901010407050d0a03f30609060001040405000603f3770908000106039401090800010421050903d502090200010404051403ea7c090400010603ad7f09080001052306032a0902000103ea00090800010603ec7e090400010417050c0603ed03090a00010404050903817d090a0001050e032e09160001060b0300090200010417050d0603d20209040001090e00000101004743433a2028292031322e322e30004c696e6b65723a204c4c442031362e302e320000000000000000000000000000000000000000000000000000000000010000000400f1ff000000000000000000000000000000000000000000000300ea2601000000000000000000000000000000000000000300ee2601000000000000000000000000000000000000000300222701000000000000000000000000001e00000000000300222701000000000000000000000000002a0000000100050008bd01000000000010000000000000005300000002000300aa880100000000004e000000000000009b0000000000030020280100000000000000000000000000a70000000100010091040100000000000c00000000000000d30000000000030064280100000000000000000000000000df000000000003008e280100000000000000000000000000eb00000002000300ca7401000000000036000000000000004501000002000300ae91010000000000080000000000000054010000020003000c950100000000002800000000000000cd010000000003007e290100000000000000000000000000d901000000000300ac290100000000000000000000000000e501000000000300d4290100000000000000000000000000f1010000020003009c7201000000000022000000000000006c02000002000300c86f010000000000d6000000000000000003000002000300be720100000000003a000000000000003903000002000300f47301000000000042000000000000007803000000000300722a010000000000000000000000000084030000000003009c2a01000000000000000000000000009003000002000300f872010000000000fc0000000000000018040000020003003a7201000000000062000000000000004b04000000000300e82b0100000000000000000000000000570400000100010056040100000000000c000000000000008204000000000300082c01000000000000000000000000008f040000010001004c040100000000000a00000000000000ba04000002000300ce710100000000006c00000000000000ed04000002000300dc90010000000000ba000000000000006e05000002000300fa8c0100000000005400000000000000af05000002000300c08f010000000000a2000000000000004c06000002000300308a0100000000005600000000000000ab060000000003009a2e0100000000000000000000000000b8060000010001009d040100000000001100000000000000e406000000000300de2e0100000000000000000000000000f106000000000300082f0100000000000000000000000000fe06000000000300982f01000000000000000000000000000b07000000000300c62f01000000000000000000000000001807000000000300ee2f010000000000000000000000000025070000000003008c3001000000000000000000000000003207000000000300b63001000000000000000000000000003f0700000200030012860100000000000e00000000000000a50700000000030064320100000000000000000000000000b20700000100010070040100000000002100000000000000bb070000020003006e7e0100000000000e00000000000000e807000002000300d09101000000000072000000000000006908000002000300fc750100000000006001000000000000a5080000020003004e8d0100000000007c01000000000000eb0800000200030098960100000000008605000000000000200900000200030000750100000000007a000000000000006109000002000300be430100000000005800000000000000b8090000020003000e430100000000005800000000000000140a000002000300664301000000000058000000000000006e0a00000200030068a30100000000008601000000000000af0a00000200030034950100000000006401000000000000e90a00000200030012450100000000005800000000000000480b000002000300b6420100000000005800000000000000a30b000002000300369f0100000000009200000000000000de0b000000000300943b0100000000000000000000000000eb0b00000100010040090100000000001c00000000000000f50b0000000003002e3c0100000000000000000000000000020c00000100010060090100000000002b000000000000002d0c000000000300363c01000000000000000000000000003a0c00000100010018020100000000002000000000000000650c000000000300403c0100000000000000000000000000720c000000000300483c01000000000000000000000000007f0c0000020003001e800100000000000e00000000000000b20c000002000300c89f010000000000a003000000000000f60c000002000300164401000000000052000000000000004f0d0000020003006a450100000000004e00000000000000a20d00000200030068440100000000005800000000000000f50d000002000300c0440100000000005200000000000000550e0000020003001e9c01000000000018030000000000008c0e00000000030014400100000000000000000000000000990e0000000003001c400100000000000000000000000000a60e000001000100b0090100000000002000000000000000d10e00000000030062410100000000000000000000000000de0e0000000003006a410100000000000000000000000000eb0e000001000100b0010100000000002000000000000000150f00000000030074410100000000000000000000000000220f0000000003007c4101000000000000000000000000002f0f0000000003008e4101000000000000000000000000003c0f00000000030096410100000000000000000000000000490f000000000300a0410100000000000000000000000000560f000000000300a8410100000000000000000000000000630f000000000300b2410100000000000000000000000000700f00000100010050070100000000002b000000000000009a0f000000000300c2410100000000000000000000000000a70f000001000100d0010100000000001c00000000000000ad0f000000000300cc410100000000000000000000000000ba0f000001000100f0010100000000002100000000000000c00f000000000300d8410100000000000000000000000000cd0f000000000300e4410100000000000000000000000000da0f000000000300f0410100000000000000000000000000000000000000030002420100000000000000000000000000e70f00000200030002420100000000000a00000000000000000000000000030002420100000000000000000000000000f90f0000020003005c77010000000000180000000000000000000000000003000c4201000000000000000000000000002e100000020003000c42010000000000080000000000000000000000000003000c42010000000000000000000000000039100000020003000268010000000000d403000000000000000000000000030014420100000000000000000000000000c41000000200030014420100000000000800000000000000000000000000030014420100000000000000000000000000d110000002000300d66b010000000000f20300000000000000000000000003001c4201000000000000000000000000005e110000020003001c420100000000004e0000000000000000000000000003001c42010000000000000000000000000000000000000003001e42010000000000000000000000000000000000000003002842010000000000000000000000000000000000000003006a4201000000000000000000000000006b110000020003006a42010000000000300000000000000000000000000003006a42010000000000000000000000000000000000000003006c42010000000000000000000000000000000000000003007242010000000000000000000000000000000000000003009a4201000000000000000000000000007d110000020003009a420100000000000e0000000000000000000000000003009a42010000000000000000000000000000000000000003009a42010000000000000000000000000000000000000003009a42010000000000000000000000000000000000000003009c42010000000000000000000000000000000000000003009c42010000000000000000000000000000000000000003009e420100000000000000000000000000b6110000020003003a800100000000000e000000000000000000000000000300a84201000000000000000000000000000000000000000300a8420100000000000000000000000000f111000002000300a8420100000000000e000000000000000000000000000300a84201000000000000000000000000000000000000000300a84201000000000000000000000000000000000000000300a84201000000000000000000000000000000000000000300aa4201000000000000000000000000000000000000000300aa4201000000000000000000000000000000000000000300ac4201000000000000000000000000000000000000000300b64201000000000000000000000000000000000000000300b64201000000000000000000000000000000000000000300b64201000000000000000000000000000000000000000300b84201000000000000000000000000000000000000000300bc420100000000000000000000000000fb11000000000300ee4201000000000000000000000000000812000000000300f642010000000000000000000000000000000000000003000e43010000000000000000000000000000000000000003000e43010000000000000000000000000000000000000003001043010000000000000000000000000000000000000003001443010000000000000000000000000015120000000003004643010000000000000000000000000022120000000003004e43010000000000000000000000000000000000000003006643010000000000000000000000000000000000000003006643010000000000000000000000000000000000000003006843010000000000000000000000000000000000000003006c4301000000000000000000000000002f120000000003009e4301000000000000000000000000003c12000000000300a64301000000000000000000000000000000000000000300be4301000000000000000000000000000000000000000300be4301000000000000000000000000000000000000000300c04301000000000000000000000000000000000000000300c44301000000000000000000000000004912000000000300f64301000000000000000000000000005612000000000300fe43010000000000000000000000000000000000000003001644010000000000000000000000000000000000000003001644010000000000000000000000000000000000000003001844010000000000000000000000000000000000000003001a4401000000000000000000000000006312000002000300428f0100000000007e00000000000000e81200000000030048440100000000000000000000000000f5120000000003005044010000000000000000000000000000000000000003006844010000000000000000000000000000000000000003006844010000000000000000000000000000000000000003006a44010000000000000000000000000000000000000003006e4401000000000000000000000000000213000000000300a04401000000000000000000000000000f13000000000300a84401000000000000000000000000000000000000000300c04401000000000000000000000000000000000000000300c04401000000000000000000000000000000000000000300c24401000000000000000000000000000000000000000300c44401000000000000000000000000001c13000002000300ca8e0100000000007800000000000000a213000000000300f2440100000000000000000000000000af13000000000300fa440100000000000000000000000000000000000000030012450100000000000000000000000000000000000000030012450100000000000000000000000000000000000000030014450100000000000000000000000000000000000000030018450100000000000000000000000000bc130000000003004a450100000000000000000000000000c9130000000003005245010000000000000000000000000000000000000003006a45010000000000000000000000000000000000000003006a45010000000000000000000000000000000000000003006c450100000000000000000000000000000000000000030070450100000000000000000000000000d61300000000030096450100000000000000000000000000e3130000000003009e4501000000000000000000000000000000000000000300b8450100000000000000000000000000f013000002000300b8450100000000009a000000000000000000000000000300b84501000000000000000000000000000000000000000300ba4501000000000000000000000000000000000000000300c24501000000000000000000000000003614000000000300d845010000000000000000000000000043140000010001003802010000000000400000000000000000000000000003005246010000000000000000000000000081140000020003005246010000000000dc00000000000000000000000000030052460100000000000000000000000000000000000000030056460100000000000000000000000000000000000000030062460100000000000000000000000000c3140000020003002e47010000000000ee1a00000000000000000000000003002e4701000000000000000000000000000715000000000400f0bb01000000000000000000000000001115000000000400f8bb01000000000000000000000000001b1500000000040000bc0100000000000000000000000000251500000000040008bc01000000000000000000000000002f1500000000040010bc0100000000000000000000000000391500000000040018bc0100000000000000000000000000431500000000040020bc01000000000000000000000000004d1500000000040028bc010000000000000000000000000000000000000003002e47010000000000000000000000000000000000000003003047010000000000000000000000000000000000000003004a4701000000000000000000000000005715000000000300ca4701000000000000000000000000006415000000000300de47010000000000000000000000000071150000000003002a4801000000000000000000000000007e150000000003003e4801000000000000000000000000008b15000000000300884801000000000000000000000000009815000000000300a2480100000000000000000000000000a515000000000300e8480100000000000000000000000000b215000000000300fe48010000000000000000000000000000000000000003001c620100000000000000000000000000bf150000020003001c62010000000000140400000000000000000000000003001c62010000000000000000000000000000000000000003001e620100000000000000000000000000000000000000030038620100000000000000000000000000011600000200030030660100000000003c000000000000003b16000000000300fe620100000000000000000000000000481600000100010060030100000000001c00000000000000511600000200030076660100000000004c000000000000008a16000002000300c2660100000000004c00000000000000d5160000020003002c800100000000000e0000000000000008170000000003007665010000000000000000000000000015170000000003008a6501000000000000000000000000002217000000000300946501000000000000000000000000002f170000000003009e6501000000000000000000000000003c17000000000300a86501000000000000000000000000004917000001000100000301000000000021000000000000005217000000000300b26501000000000000000000000000005f17000001000100300301000000000024000000000000006817000000000300c06501000000000000000000000000007517000000000300ca6501000000000000000000000000008217000001000100d00201000000000021000000000000008b17000000000300d46501000000000000000000000000009817000000000300de650100000000000000000000000000a517000000000300e8650100000000000000000000000000b217000001000100a0020100000000002300000000000000bb17000000000300f6650100000000000000000000000000c817000001000100a0030100000000001000000000000000f317000000000300106601000000000000000000000000000018000001000100e80301000000000010000000000000002b180000020003006c660100000000000a000000000000006118000000000300226601000000000000000000000000000000000000000300306601000000000000000000000000000000000000000300306601000000000000000000000000006e18000000000300486601000000000000000000000000007b180000000003005666010000000000000000000000000000000000000003006c66010000000000000000000000000000000000000003006c66010000000000000000000000000000000000000003007666010000000000000000000000000000000000000003007666010000000000000000000000000088180000000003009466010000000000000000000000000095180000000003009e660100000000000000000000000000a218000000000300ac6601000000000000000000000000000000000000000300c26601000000000000000000000000000000000000000300c2660100000000000000000000000000af18000000000300e2660100000000000000000000000000bc18000000000300ec660100000000000000000000000000c91800000000030002670100000000000000000000000000d618000001000100f8030100000000000d0000000000000000000000000003000e67010000000000000000000000000001190000020003000e67010000000000f40000000000000000000000000003000e6701000000000000000000000000004019000000000300da6701000000000000000000000000004d19000000000300ee6701000000000000000000000000005a19000000000300f867010000000000000000000000000000000000000003000268010000000000000000000000000000000000000003000268010000000000000000000000000000000000000003000468010000000000000000000000000000000000000003001c680100000000000000000000000000671900000000030022680100000000000000000000000000741900000100050060bc010000000000a80000000000000098190000000003002e680100000000000000000000000000a519000000000300d8690100000000000000000000000000b3190000000003001a6a0100000000000000000000000000c1190000000003004a6b0100000000000000000000000000cf19000000000300546b0100000000000000000000000000dd19000000000300626b0100000000000000000000000000eb19000000000300766b0100000000000000000000000000f919000000000300806b0100000000000000000000000000061a000000000300946b0100000000000000000000000000131a0000000003009c6b0100000000000000000000000000211a000001000100780201000000000020000000000000004b1a000000000300a66b0100000000000000000000000000581a000000000300ae6b0100000000000000000000000000651a000000000300b86b0100000000000000000000000000731a000000000300c06b01000000000000000000000000000000000000000300d66b01000000000000000000000000000000000000000300d66b01000000000000000000000000000000000000000300d86b01000000000000000000000000000000000000000300f26b0100000000000000000000000000811a000000000300f26b01000000000000000000000000008f1a000000000300106c01000000000000000000000000009d1a0000000003005c6c0100000000000000000000000000ab1a000000000300046d0100000000000000000000000000b91a000000000300546f0100000000000000000000000000c71a0000000003005e6f0100000000000000000000000000d51a0000000003006c6f0100000000000000000000000000e31a000000000300806f0100000000000000000000000000f11a000000000300986f0100000000000000000000000000ff1a000000000300a06f01000000000000000000000000000d1b000000000300aa6f01000000000000000000000000001b1b000000000300b26f01000000000000000000000000000000000000000300c86f01000000000000000000000000000000000000000300c86f01000000000000000000000000000000000000000300ca6f01000000000000000000000000000000000000000300d86f0100000000000000000000000000291b0000020003009e700100000000005200000000000000711b000002000300f0700100000000003400000000000000cb1b0000000003007c700100000000000000000000000000d91b0000010001001004010000000000190000000000000000000000000003009e70010000000000000000000000000000000000000003009e7001000000000000000000000000000000000000000300a07001000000000000000000000000000000000000000300a6700100000000000000000000000000e21b000002000300a6910100000000000800000000000000ef1b000002000300c6910100000000000a000000000000000000000000000300f07001000000000000000000000000000000000000000300f07001000000000000000000000000000000000000000300f27001000000000000000000000000000000000000000300f47001000000000000000000000000000a1c0000020003002471010000000000740000000000000000000000000003002471010000000000000000000000000000000000000003002471010000000000000000000000000000000000000003002671010000000000000000000000000000000000000003002c710100000000000000000000000000551c00000200030018880100000000006200000000000000000000000000030098710100000000000000000000000000881c0000020003009871010000000000360000000000000000000000000003009871010000000000000000000000000000000000000003009a71010000000000000000000000000000000000000003009c7101000000000000000000000000000000000000000300ce7101000000000000000000000000000000000000000300ce7101000000000000000000000000000000000000000300d07101000000000000000000000000000000000000000300dc71010000000000000000000000000000000000000003003a72010000000000000000000000000000000000000003003a72010000000000000000000000000000000000000003003c72010000000000000000000000000000000000000003004872010000000000000000000000000000000000000003009c72010000000000000000000000000000000000000003009c7201000000000000000000000000000000000000000300be7201000000000000000000000000000000000000000300be7201000000000000000000000000000000000000000300c07201000000000000000000000000000000000000000300c67201000000000000000000000000000000000000000300f87201000000000000000000000000000000000000000300f87201000000000000000000000000000000000000000300fa720100000000000000000000000000000000000000030008730100000000000000000000000000d51c00000000030024730100000000000000000000000000e31c00000100010062040100000000000b000000000000000f1d000000000300807301000000000000000000000000001d1d000000000300da7301000000000000000000000000000000000000000300f47301000000000000000000000000000000000000000300f47301000000000000000000000000000000000000000300367401000000000000000000000000002b1d0000020003003674010000000000920000000000000000000000000003003674010000000000000000000000000000000000000003003874010000000000000000000000000000000000000003003a740100000000000000000000000000861d0000000003003e740100000000000000000000000000941d000000000100600101000000000000000000000000009e1d0000000003004c740100000000000000000000000000a71d00000000030052740100000000000000000000000000b51d0000010001002b050100000000000f00000000000000e01d0000000003005e740100000000000000000000000000e91d00000000030064740100000000000000000000000000f71d00000100010020050100000000000b00000000000000221e000000000300707401000000000000000000000000002b1e00000000030074740100000000000000000000000000391e000001000100f0040100000000000f00000000000000641e0000000003007c740100000000000000000000000000721e000001000100000501000000000020000000000000009d1e00000000030088740100000000000000000000000000a61e0000000003008e740100000000000000000000000000b41e0000000003009e740100000000000000000000000000bd1e000000000300a2740100000000000000000000000000cb1e000001000100ae040100000000000700000000000000f61e000000000300aa740100000000000000000000000000041f000001000100b80401000000000020000000000000002f1f0000020003007a8501000000000098000000000000000000000000000300c8740100000000000000000000000000751f000002000300c87401000000000002000000000000000000000000000300c87401000000000000000000000000000000000000000300ca7401000000000000000000000000000000000000000300ca74010000000000000000000000000000000000000003000075010000000000000000000000000000000000000003000075010000000000000000000000000000000000000003000275010000000000000000000000000000000000000003000675010000000000000000000000000000000000000003007a750100000000000000000000000000b41f0000020003007a75010000000000820000000000000000000000000003007a75010000000000000000000000000000000000000003007c7501000000000000000000000000000000000000000300807501000000000000000000000000000000000000000300fc7501000000000000000000000000000000000000000300fc75010000000000000000000000000000000000000003000076010000000000000000000000000000000000000003002476010000000000000000000000000000000000000003005c77010000000000000000000000000000000000000003005c770100000000000000000000000000000000000000030074770100000000000000000000000000f51f0000020003007477010000000000040000000000000000000000000003007477010000000000000000000000000000000000000003007477010000000000000000000000000000000000000003007477010000000000000000000000000000000000000003007477010000000000000000000000000000000000000003007677010000000000000000000000000000000000000003007677010000000000000000000000000000000000000003007877010000000000000000000000000000000000000003007877010000000000000000000000000000000000000003007877010000000000000000000000000030200000020003007877010000000000020000000000000000000000000003007877010000000000000000000000000000000000000003007877010000000000000000000000000000000000000003007877010000000000000000000000000000000000000003007877010000000000000000000000000000000000000003007a77010000000000000000000000000000000000000003007a770100000000000000000000000000ba2000000000040030bc0100000000000000000000000000c4200000020003007a77010000000000420100000000000000000000000003007a77010000000000000000000000000000000000000003007a77010000000000000000000000000000000000000003007a77010000000000000000000000000000000000000003007c77010000000000000000000000000000000000000003007e770100000000000000000000000000000000000000030080770100000000000000000000000000f5200000000003008c77010000000000000000000000000003210000010001009e05010000000000c80000000000000000000000000003009877010000000000000000000000000000000000000003009c7701000000000000000000000000002f21000000000300a07701000000000000000000000000000000000000000300c07701000000000000000000000000000000000000000300c27701000000000000000000000000000000000000000300d07701000000000000000000000000000000000000000300ea7701000000000000000000000000000000000000000300ea7701000000000000000000000000000000000000000300ec7701000000000000000000000000000000000000000300ec7701000000000000000000000000000000000000000300f07701000000000000000000000000000000000000000300f07701000000000000000000000000000000000000000300f47701000000000000000000000000000000000000000300f47701000000000000000000000000000000000000000300fc7701000000000000000000000000000000000000000300fc7701000000000000000000000000000000000000000300fe7701000000000000000000000000000000000000000300fe77010000000000000000000000000000000000000003000678010000000000000000000000000000000000000003000678010000000000000000000000000000000000000003000878010000000000000000000000000000000000000003000878010000000000000000000000000000000000000003000c78010000000000000000000000000000000000000003000c78010000000000000000000000000000000000000003001478010000000000000000000000000000000000000003001478010000000000000000000000000000000000000003001a78010000000000000000000000000000000000000003001e78010000000000000000000000000000000000000003002278010000000000000000000000000000000000000003003e78010000000000000000000000000000000000000003004278010000000000000000000000000000000000000003004478010000000000000000000000000000000000000003004478010000000000000000000000000000000000000003004678010000000000000000000000000000000000000003004678010000000000000000000000000000000000000003005278010000000000000000000000000000000000000003005278010000000000000000000000000000000000000003005478010000000000000000000000000000000000000003005478010000000000000000000000000000000000000003005e78010000000000000000000000000000000000000003005e78010000000000000000000000000000000000000003006078010000000000000000000000000000000000000003006478010000000000000000000000000000000000000003006c78010000000000000000000000000000000000000003006c78010000000000000000000000000000000000000003006e78010000000000000000000000000000000000000003006e78010000000000000000000000000000000000000003007878010000000000000000000000000000000000000003007a78010000000000000000000000000000000000000003007e78010000000000000000000000000000000000000003007e78010000000000000000000000000000000000000003008078010000000000000000000000000000000000000003008078010000000000000000000000000000000000000003008c78010000000000000000000000000000000000000003008c78010000000000000000000000000000000000000003008e78010000000000000000000000000000000000000003008e78010000000000000000000000000000000000000003009678010000000000000000000000000000000000000003009678010000000000000000000000000000000000000003009a78010000000000000000000000000000000000000003009a7801000000000000000000000000000000000000000300a07801000000000000000000000000000000000000000300a07801000000000000000000000000003d21000000000300a27801000000000000000000000000004b21000001000100600901000000000000000000000000000000000000000300a27801000000000000000000000000007621000002000300bc78010000000000e4010000000000000000000000000300b67801000000000000000000000000000000000000000300b87801000000000000000000000000000000000000000300bc7801000000000000000000000000000000000000000300bc7801000000000000000000000000000000000000000300bc7801000000000000000000000000000000000000000300bc7801000000000000000000000000000000000000000300bc7801000000000000000000000000000000000000000300be7801000000000000000000000000000000000000000300d87801000000000000000000000000000000000000000300da7801000000000000000000000000000000000000000300da7801000000000000000000000000000000000000000300e67801000000000000000000000000000000000000000300e67801000000000000000000000000000000000000000300f27801000000000000000000000000000000000000000300f67801000000000000000000000000000000000000000300f67801000000000000000000000000000000000000000300fa7801000000000000000000000000000000000000000300fa7801000000000000000000000000000000000000000300fc7801000000000000000000000000000000000000000300fe78010000000000000000000000000000000000000003000079010000000000000000000000000000000000000003000279010000000000000000000000000000000000000003000679010000000000000000000000000000000000000003000879010000000000000000000000000000000000000003000879010000000000000000000000000000000000000003000c79010000000000000000000000000000000000000003000c79010000000000000000000000000000000000000003001079010000000000000000000000000000000000000003001479010000000000000000000000000000000000000003001479010000000000000000000000000000000000000003001679010000000000000000000000000000000000000003001679010000000000000000000000000000000000000003001e79010000000000000000000000000000000000000003001e79010000000000000000000000000000000000000003002079010000000000000000000000000000000000000003002079010000000000000000000000000000000000000003002279010000000000000000000000000000000000000003002279010000000000000000000000000000000000000003002479010000000000000000000000000000000000000003002479010000000000000000000000000000000000000003002679010000000000000000000000000000000000000003002879010000000000000000000000000000000000000003002a79010000000000000000000000000000000000000003002e79010000000000000000000000000000000000000003003279010000000000000000000000000000000000000003003279010000000000000000000000000000000000000003003479010000000000000000000000000000000000000003003479010000000000000000000000000000000000000003003679010000000000000000000000000000000000000003003679010000000000000000000000000000000000000003003c79010000000000000000000000000000000000000003003c790100000000000000000000000000000000000000030040790100000000000000000000000000000000000000030040790100000000000000000000000000000000000000030046790100000000000000000000000000000000000000030046790100000000000000000000000000af21000002000300a07a01000000000056000000000000000000000000000300667901000000000000000000000000000000000000000300827901000000000000000000000000000000000000000300867901000000000000000000000000000000000000000300ac7901000000000000000000000000000000000000000300ac7901000000000000000000000000000000000000000300b27901000000000000000000000000000000000000000300b27901000000000000000000000000000000000000000300b67901000000000000000000000000000000000000000300b67901000000000000000000000000000000000000000300c07901000000000000000000000000000000000000000300c07901000000000000000000000000000000000000000300c47901000000000000000000000000000000000000000300c47901000000000000000000000000000000000000000300c87901000000000000000000000000000000000000000300c87901000000000000000000000000000000000000000300dc7901000000000000000000000000000000000000000300de7901000000000000000000000000000000000000000300de7901000000000000000000000000000000000000000300e47901000000000000000000000000000000000000000300e47901000000000000000000000000000000000000000300e87901000000000000000000000000000000000000000300e87901000000000000000000000000000000000000000300f87901000000000000000000000000000000000000000300f87901000000000000000000000000000000000000000300fa7901000000000000000000000000000000000000000300fa7901000000000000000000000000000000000000000300fe7901000000000000000000000000000000000000000300027a01000000000000000000000000000000000000000300047a010000000000000000000000000000000000000003000a7a01000000000000000000000000000000000000000300167a010000000000000000000000000000000000000003001a7a010000000000000000000000000000000000000003001a7a010000000000000000000000000000000000000003001c7a010000000000000000000000000000000000000003001c7a010000000000000000000000000000000000000003001e7a010000000000000000000000000000000000000003001e7a010000000000000000000000000000000000000003002a7a010000000000000000000000000000000000000003002a7a01000000000000000000000000000000000000000300347a01000000000000000000000000000000000000000300387a010000000000000000000000000000000000000003004c7a010000000000000000000000000000000000000003005a7a010000000000000000000000000000000000000003005a7a01000000000000000000000000000000000000000300627a01000000000000000000000000000000000000000300627a010000000000000000000000000000000000000003006a7a010000000000000000000000000000000000000003006a7a010000000000000000000000000000000000000003007a7a010000000000000000000000000000000000000003007a7a010000000000000000000000000000000000000003008a7a010000000000000000000000000000000000000003008c7a01000000000000000000000000000000000000000300907a01000000000000000000000000000000000000000300987a010000000000000000000000000000000000000003009a7a010000000000000000000000000000000000000003009a7a01000000000000000000000000000000000000000300a07a01000000000000000000000000000000000000000300a07a01000000000000000000000000000000000000000300a07a01000000000000000000000000000000000000000300a07a01000000000000000000000000000000000000000300a07a01000000000000000000000000000000000000000300a07a01000000000000000000000000000000000000000300a27a01000000000000000000000000000000000000000300ac7a01000000000000000000000000000000000000000300bc7a01000000000000000000000000000000000000000300c07a01000000000000000000000000000000000000000300ce7a01000000000000000000000000000000000000000300d07a01000000000000000000000000000000000000000300e27a01000000000000000000000000000000000000000300e67a01000000000000000000000000000000000000000300e87a01000000000000000000000000000000000000000300f27a01000000000000000000000000000000000000000300f67a01000000000000000000000000000000000000000300f67a0100000000000000000000000000f62100000000040038bc0100000000000000000000000000002200000000040040bc01000000000000000000000000000a22000002000300f67a01000000000078030000000000000000000000000300f67a01000000000000000000000000000000000000000300f67a01000000000000000000000000000000000000000300f67a01000000000000000000000000000000000000000300f87a01000000000000000000000000000000000000000300f87a01000000000000000000000000000000000000000300f87a010000000000000000000000000000000000000003000a7b010000000000000000000000000000000000000003000e7b010000000000000000000000000000000000000003000e7b01000000000000000000000000000000000000000300107b01000000000000000000000000000000000000000300107b01000000000000000000000000000000000000000300187b01000000000000000000000000000000000000000300187b010000000000000000000000000000000000000003001c7b01000000000000000000000000000000000000000300207b01000000000000000000000000000000000000000300247b01000000000000000000000000000000000000000300247b01000000000000000000000000000000000000000300287b01000000000000000000000000000000000000000300287b010000000000000000000000000000000000000003003a7b010000000000000000000000000000000000000003003a7b010000000000000000000000000000000000000003003e7b010000000000000000000000000000000000000003003e7b01000000000000000000000000000000000000000300407b01000000000000000000000000000000000000000300447b01000000000000000000000000000000000000000300447b01000000000000000000000000000000000000000300487b01000000000000000000000000000000000000000300487b010000000000000000000000000000000000000003004a7b010000000000000000000000000000000000000003004a7b010000000000000000000000000000000000000003004c7b010000000000000000000000000000000000000003004c7b01000000000000000000000000000000000000000300507b01000000000000000000000000000000000000000300507b01000000000000000000000000000000000000000300587b010000000000000000000000000000000000000003005c7b01000000000000000000000000000000000000000300607b01000000000000000000000000000000000000000300607b01000000000000000000000000000000000000000300647b01000000000000000000000000000000000000000300647b01000000000000000000000000000000000000000300687b01000000000000000000000000000000000000000300687b010000000000000000000000000000000000000003006c7b01000000000000000000000000000000000000000300707b01000000000000000000000000000000000000000300707b01000000000000000000000000000000000000000300727b01000000000000000000000000000000000000000300767b010000000000000000000000000000000000000003007a7b010000000000000000000000000000000000000003007a7b010000000000000000000000000000000000000003007e7b01000000000000000000000000000000000000000300827b01000000000000000000000000000000000000000300867b01000000000000000000000000000000000000000300867b01000000000000000000000000000000000000000300887b010000000000000000000000000000000000000003008c7b01000000000000000000000000000000000000000300907b01000000000000000000000000000000000000000300907b01000000000000000000000000000000000000000300927b01000000000000000000000000000000000000000300927b01000000000000000000000000000000000000000300967b01000000000000000000000000000000000000000300967b01000000000000000000000000000000000000000300b47b01000000000000000000000000000000000000000300b47b01000000000000000000000000000000000000000300b87b01000000000000000000000000000000000000000300b87b01000000000000000000000000000000000000000300bc7b01000000000000000000000000000000000000000300c07b01000000000000000000000000000000000000000300c87b01000000000000000000000000000000000000000300cc7b01000000000000000000000000000000000000000300d07b01000000000000000000000000000000000000000300d47b01000000000000000000000000000000000000000300d87b01000000000000000000000000000000000000000300dc7b01000000000000000000000000000000000000000300dc7b01000000000000000000000000000000000000000300e07b01000000000000000000000000000000000000000300e07b01000000000000000000000000000000000000000300e47b01000000000000000000000000000000000000000300e47b01000000000000000000000000000000000000000300e87b01000000000000000000000000000000000000000300ec7b01000000000000000000000000000000000000000300ec7b01000000000000000000000000000000000000000300f27b01000000000000000000000000000000000000000300f67b01000000000000000000000000000000000000000300f87b01000000000000000000000000000000000000000300f87b01000000000000000000000000000000000000000300fe7b01000000000000000000000000000000000000000300fe7b01000000000000000000000000000000000000000300027c01000000000000000000000000000000000000000300027c01000000000000000000000000000000000000000300047c01000000000000000000000000000000000000000300087c01000000000000000000000000000000000000000300087c010000000000000000000000000000000000000003000c7c010000000000000000000000000000000000000003000c7c01000000000000000000000000000000000000000300147c01000000000000000000000000000000000000000300147c01000000000000000000000000000000000000000300187c01000000000000000000000000000000000000000300187c010000000000000000000000000000000000000003001a7c010000000000000000000000000000000000000003001a7c010000000000000000000000000000000000000003001e7c010000000000000000000000000000000000000003001e7c01000000000000000000000000000000000000000300227c01000000000000000000000000000000000000000300227c01000000000000000000000000000000000000000300247c01000000000000000000000000000000000000000300247c01000000000000000000000000000000000000000300267c01000000000000000000000000000000000000000300267c010000000000000000000000000000000000000003002a7c010000000000000000000000000000000000000003002e7c01000000000000000000000000000000000000000300367c01000000000000000000000000000000000000000300367c010000000000000000000000000000000000000003003a7c010000000000000000000000000000000000000003003c7c010000000000000000000000000000000000000003003c7c01000000000000000000000000000000000000000300407c01000000000000000000000000000000000000000300407c01000000000000000000000000000000000000000300447c01000000000000000000000000000000000000000300487c01000000000000000000000000000000000000000300487c010000000000000000000000000000000000000003004a7c010000000000000000000000000000000000000003004a7c01000000000000000000000000000000000000000300527c01000000000000000000000000000000000000000300527c01000000000000000000000000000000000000000300547c01000000000000000000000000000000000000000300547c01000000000000000000000000000000000000000300567c01000000000000000000000000000000000000000300567c010000000000000000000000000000000000000003005a7c010000000000000000000000000000000000000003005a7c01000000000000000000000000000000000000000300607c01000000000000000000000000000000000000000300607c01000000000000000000000000000000000000000300687c01000000000000000000000000000000000000000300687c010000000000000000000000000000000000000003006e7c010000000000000000000000000000000000000003006e7c01000000000000000000000000000000000000000300727c01000000000000000000000000000000000000000300727c01000000000000000000000000000000000000000300747c01000000000000000000000000000000000000000300787c01000000000000000000000000000000000000000300787c010000000000000000000000000000000000000003007a7c010000000000000000000000000000000000000003007a7c01000000000000000000000000000000000000000300827c01000000000000000000000000000000000000000300827c01000000000000000000000000000000000000000300847c01000000000000000000000000000000000000000300847c01000000000000000000000000000000000000000300867c01000000000000000000000000000000000000000300867c01000000000000000000000000000000000000000300887c01000000000000000000000000000000000000000300887c010000000000000000000000000000000000000003008a7c010000000000000000000000000000000000000003008a7c010000000000000000000000000000000000000003008c7c010000000000000000000000000000000000000003008c7c01000000000000000000000000000000000000000300927c01000000000000000000000000000000000000000300967c01000000000000000000000000000000000000000300967c01000000000000000000000000000000000000000300987c01000000000000000000000000000000000000000300987c01000000000000000000000000000000000000000300a07c01000000000000000000000000000000000000000300a07c01000000000000000000000000000000000000000300a27c01000000000000000000000000000000000000000300a27c01000000000000000000000000000000000000000300a47c01000000000000000000000000000000000000000300a47c01000000000000000000000000000000000000000300a67c01000000000000000000000000000000000000000300a67c01000000000000000000000000003922000000000300aa7c01000000000000000000000000004722000000000300b27c01000000000000000000000000000000000000000300c87c01000000000000000000000000000000000000000300ce7c01000000000000000000000000000000000000000300dc7c01000000000000000000000000000000000000000300dc7c01000000000000000000000000000000000000000300e07c01000000000000000000000000000000000000000300e27c01000000000000000000000000000000000000000300e67c01000000000000000000000000000000000000000300e87c01000000000000000000000000000000000000000300e87c01000000000000000000000000000000000000000300ec7c01000000000000000000000000000000000000000300ec7c01000000000000000000000000000000000000000300ee7c01000000000000000000000000000000000000000300ee7c01000000000000000000000000000000000000000300f07c01000000000000000000000000000000000000000300f27c01000000000000000000000000000000000000000300f27c01000000000000000000000000000000000000000300f47c01000000000000000000000000000000000000000300fe7c01000000000000000000000000000000000000000300027d01000000000000000000000000000000000000000300067d01000000000000000000000000000000000000000300067d010000000000000000000000000000000000000003000a7d010000000000000000000000000000000000000003000a7d01000000000000000000000000000000000000000300107d01000000000000000000000000000000000000000300107d01000000000000000000000000000000000000000300127d01000000000000000000000000000000000000000300127d01000000000000000000000000000000000000000300167d01000000000000000000000000000000000000000300187d010000000000000000000000000000000000000003001a7d010000000000000000000000000000000000000003001a7d010000000000000000000000000000000000000003001e7d01000000000000000000000000000000000000000300207d01000000000000000000000000000000000000000300227d01000000000000000000000000000000000000000300227d01000000000000000000000000000000000000000300247d01000000000000000000000000000000000000000300247d01000000000000000000000000000000000000000300287d01000000000000000000000000000000000000000300287d010000000000000000000000000000000000000003002a7d010000000000000000000000000000000000000003002a7d010000000000000000000000000000000000000003002e7d01000000000000000000000000000000000000000300307d01000000000000000000000000000000000000000300307d01000000000000000000000000000000000000000300327d01000000000000000000000000000000000000000300327d01000000000000000000000000000000000000000300347d01000000000000000000000000000000000000000300387d010000000000000000000000000000000000000003003c7d010000000000000000000000000000000000000003003e7d01000000000000000000000000000000000000000300407d01000000000000000000000000000000000000000300427d01000000000000000000000000000000000000000300427d01000000000000000000000000000000000000000300447d01000000000000000000000000000000000000000300447d01000000000000000000000000000000000000000300467d01000000000000000000000000000000000000000300467d010000000000000000000000000000000000000003004a7d010000000000000000000000000000000000000003004a7d010000000000000000000000000000000000000003004e7d01000000000000000000000000000000000000000300507d01000000000000000000000000000000000000000300527d01000000000000000000000000000000000000000300567d01000000000000000000000000000000000000000300567d010000000000000000000000000000000000000003005a7d010000000000000000000000000000000000000003005a7d010000000000000000000000000000000000000003005c7d010000000000000000000000000000000000000003005c7d01000000000000000000000000000000000000000300627d01000000000000000000000000000000000000000300627d01000000000000000000000000000000000000000300667d010000000000000000000000000000000000000003006a7d010000000000000000000000000000000000000003006e7d01000000000000000000000000000000000000000300747d010000000000000000000000000000000000000003007a7d010000000000000000000000000000000000000003007a7d010000000000000000000000000000000000000003007c7d010000000000000000000000000000000000000003007c7d010000000000000000000000000000000000000003007e7d010000000000000000000000000000000000000003007e7d01000000000000000000000000000000000000000300827d01000000000000000000000000000000000000000300847d01000000000000000000000000000000000000000300867d010000000000000000000000000000000000000003008a7d010000000000000000000000000000000000000003008a7d010000000000000000000000000000000000000003008c7d010000000000000000000000000000000000000003008c7d010000000000000000000000000000000000000003008e7d010000000000000000000000000000000000000003008e7d01000000000000000000000000000000000000000300927d01000000000000000000000000000000000000000300927d01000000000000000000000000000000000000000300947d01000000000000000000000000000000000000000300947d01000000000000000000000000000000000000000300987d010000000000000000000000000000000000000003009a7d010000000000000000000000000000000000000003009e7d01000000000000000000000000000000000000000300a07d01000000000000000000000000000000000000000300a07d01000000000000000000000000000000000000000300a47d01000000000000000000000000000000000000000300a47d01000000000000000000000000000000000000000300a67d01000000000000000000000000000000000000000300a67d01000000000000000000000000000000000000000300a87d01000000000000000000000000000000000000000300a87d01000000000000000000000000000000000000000300ac7d01000000000000000000000000000000000000000300ac7d01000000000000000000000000000000000000000300b27d01000000000000000000000000000000000000000300b27d01000000000000000000000000000000000000000300b67d01000000000000000000000000000000000000000300b67d01000000000000000000000000000000000000000300bc7d01000000000000000000000000000000000000000300bc7d01000000000000000000000000000000000000000300e27d01000000000000000000000000000000000000000300e27d01000000000000000000000000000000000000000300e67d01000000000000000000000000000000000000000300ea7d01000000000000000000000000000000000000000300ec7d01000000000000000000000000000000000000000300f27d01000000000000000000000000000000000000000300007e01000000000000000000000000000000000000000300047e01000000000000000000000000000000000000000300047e01000000000000000000000000000000000000000300067e01000000000000000000000000000000000000000300067e01000000000000000000000000000000000000000300087e01000000000000000000000000000000000000000300087e01000000000000000000000000000000000000000300147e01000000000000000000000000000000000000000300147e010000000000000000000000000000000000000003001e7e01000000000000000000000000000000000000000300227e01000000000000000000000000000000000000000300307e01000000000000000000000000000000000000000300307e01000000000000000000000000000000000000000300387e01000000000000000000000000000000000000000300387e010000000000000000000000000000000000000003003c7e010000000000000000000000000000000000000003003c7e01000000000000000000000000000000000000000300407e01000000000000000000000000000000000000000300407e01000000000000000000000000000000000000000300507e01000000000000000000000000000000000000000300527e01000000000000000000000000000000000000000300527e01000000000000000000000000000000000000000300567e01000000000000000000000000000000000000000300567e010000000000000000000000000000000000000003006a7e010000000000000000000000000000000000000003006e7e010000000000000000000000000000000000000003006e7e010000000000000000000000000000000000000003006e7e010000000000000000000000000000000000000003006e7e010000000000000000000000000000000000000003006e7e01000000000000000000000000000000000000000300707e01000000000000000000000000000000000000000300707e01000000000000000000000000000000000000000300727e010000000000000000000000000000000000000003007c7e010000000000000000000000000000000000000003007c7e010000000000000000000000000055220000020003007c7e0100000000007e0100000000000000000000000003007c7e010000000000000000000000000000000000000003007c7e010000000000000000000000000000000000000003007c7e010000000000000000000000000000000000000003007e7e010000000000000000000000000000000000000003008e7e01000000000000000000000000000000000000000300947e01000000000000000000000000000000000000000300947e010000000000000000000000000000000000000003009c7e010000000000000000000000000000000000000003009c7e01000000000000000000000000000000000000000300a07e01000000000000000000000000000000000000000300a07e01000000000000000000000000000000000000000300a87e01000000000000000000000000000000000000000300a87e01000000000000000000000000000000000000000300aa7e01000000000000000000000000000000000000000300ae7e01000000000000000000000000000000000000000300ae7e01000000000000000000000000000000000000000300b27e01000000000000000000000000000000000000000300b67e01000000000000000000000000007c22000000000300d07e01000000000000000000000000000000000000000300d87e01000000000000000000000000000000000000000300d87e01000000000000000000000000000000000000000300da7e01000000000000000000000000000000000000000300dc7e01000000000000000000000000000000000000000300e07e01000000000000000000000000000000000000000300e47e01000000000000000000000000000000000000000300ea7e01000000000000000000000000000000000000000300ea7e01000000000000000000000000000000000000000300ec7e01000000000000000000000000000000000000000300ee7e01000000000000000000000000000000000000000300f27e01000000000000000000000000000000000000000300f67e01000000000000000000000000000000000000000300f87e01000000000000000000000000000000000000000300f87e01000000000000000000000000000000000000000300fc7e01000000000000000000000000000000000000000300fc7e01000000000000000000000000000000000000000300fe7e01000000000000000000000000000000000000000300047f01000000000000000000000000000000000000000300047f010000000000000000000000000000000000000003000a7f010000000000000000000000000000000000000003000a7f01000000000000000000000000000000000000000300147f01000000000000000000000000000000000000000300187f010000000000000000000000000000000000000003001a7f010000000000000000000000000000000000000003001c7f010000000000000000000000000000000000000003001c7f010000000000000000000000000000000000000003001e7f01000000000000000000000000000000000000000300227f010000000000000000000000000000000000000003002a7f010000000000000000000000000000000000000003002a7f01000000000000000000000000000000000000000300307f01000000000000000000000000000000000000000300307f010000000000000000000000000000000000000003003a7f010000000000000000000000000000000000000003003e7f01000000000000000000000000000000000000000300407f01000000000000000000000000000000000000000300427f01000000000000000000000000000000000000000300427f01000000000000000000000000000000000000000300447f01000000000000000000000000000000000000000300487f010000000000000000000000000000000000000003004a7f010000000000000000000000000000000000000003004a7f010000000000000000000000000000000000000003004e7f010000000000000000000000000000000000000003004e7f01000000000000000000000000000000000000000300507f01000000000000000000000000000000000000000300527f01000000000000000000000000000000000000000300567f01000000000000000000000000000000000000000300567f01000000000000000000000000000000000000000300587f01000000000000000000000000000000000000000300587f01000000000000000000000000000000000000000300687f01000000000000000000000000000000000000000300687f010000000000000000000000000000000000000003006c7f010000000000000000000000000000000000000003006c7f01000000000000000000000000000000000000000300707f01000000000000000000000000000000000000000300787f010000000000000000000000000000000000000003008a7f010000000000000000000000000000000000000003008a7f010000000000000000000000000000000000000003008c7f010000000000000000000000000000000000000003008e7f01000000000000000000000000000000000000000300927f01000000000000000000000000000000000000000300967f010000000000000000000000000000000000000003009c7f010000000000000000000000000000000000000003009c7f010000000000000000000000000000000000000003009e7f01000000000000000000000000000000000000000300a27f01000000000000000000000000000000000000000300a67f01000000000000000000000000000000000000000300a67f01000000000000000000000000000000000000000300a87f01000000000000000000000000000000000000000300a87f01000000000000000000000000000000000000000300b27f01000000000000000000000000000000000000000300b27f01000000000000000000000000000000000000000300b67f01000000000000000000000000000000000000000300b67f01000000000000000000000000000000000000000300bc7f01000000000000000000000000000000000000000300bc7f01000000000000000000000000000000000000000300be7f01000000000000000000000000000000000000000300c27f01000000000000000000000000000000000000000300c27f01000000000000000000000000000000000000000300c67f01000000000000000000000000000000000000000300c67f01000000000000000000000000000000000000000300ca7f01000000000000000000000000000000000000000300ca7f01000000000000000000000000000000000000000300ce7f01000000000000000000000000000000000000000300ce7f01000000000000000000000000000000000000000300d27f01000000000000000000000000000000000000000300da7f01000000000000000000000000000000000000000300e07f01000000000000000000000000000000000000000300e67f01000000000000000000000000000000000000000300f67f01000000000000000000000000000000000000000300fa7f01000000000000000000000000000000000000000300fa7f01000000000000000000000000008a22000002000300fa7f01000000000012000000000000000000000000000300fa7f01000000000000000000000000000000000000000300fa7f01000000000000000000000000000000000000000300fa7f01000000000000000000000000000000000000000300fa7f0100000000000000000000000000e42200000000030000800100000000000000000000000000f2220000010001003b050100000000000b0000000000000000000000000003000c80010000000000000000000000000000000000000003000c80010000000000000000000000000000000000000003000c8001000000000000000000000000001e230000020003000c80010000000000120000000000000000000000000003000c80010000000000000000000000000000000000000003000c80010000000000000000000000000000000000000003000c80010000000000000000000000000000000000000003000c8001000000000000000000000000007b2300000000030012800100000000000000000000000000892300000100010046050100000000000e0000000000000000000000000003001e80010000000000000000000000000000000000000003001e80010000000000000000000000000000000000000003001e80010000000000000000000000000000000000000003001e80010000000000000000000000000000000000000003001e80010000000000000000000000000000000000000003001e80010000000000000000000000000000000000000003002080010000000000000000000000000000000000000003002080010000000000000000000000000000000000000003002280010000000000000000000000000000000000000003002c80010000000000000000000000000000000000000003002c80010000000000000000000000000000000000000003002c80010000000000000000000000000000000000000003002c80010000000000000000000000000000000000000003002c80010000000000000000000000000000000000000003002e80010000000000000000000000000000000000000003002e80010000000000000000000000000000000000000003002e80010000000000000000000000000000000000000003003080010000000000000000000000000000000000000003003a80010000000000000000000000000000000000000003003a80010000000000000000000000000000000000000003003a80010000000000000000000000000000000000000003003a80010000000000000000000000000000000000000003003a80010000000000000000000000000000000000000003003a80010000000000000000000000000000000000000003003c80010000000000000000000000000000000000000003003c80010000000000000000000000000000000000000003003e800100000000000000000000000000000000000000030048800100000000000000000000000000000000000000030048800100000000000000000000000000b5230000020003004880010000000000700000000000000000000000000003004880010000000000000000000000000000000000000003004880010000000000000000000000000000000000000003004880010000000000000000000000000000000000000003004a80010000000000000000000000000000000000000003004c80010000000000000000000000000000000000000003004e80010000000000000000000000000000000000000003004e80010000000000000000000000000000000000000003005680010000000000000000000000000000000000000003005680010000000000000000000000000000000000000003005e80010000000000000000000000000000000000000003005e80010000000000000000000000000000000000000003006080010000000000000000000000000000000000000003006080010000000000000000000000000000000000000003006480010000000000000000000000000000000000000003006480010000000000000000000000000000000000000003006c80010000000000000000000000000000000000000003006e80010000000000000000000000000000000000000003006e80010000000000000000000000000000000000000003007680010000000000000000000000000000000000000003007680010000000000000000000000000000000000000003007a80010000000000000000000000000000000000000003007a80010000000000000000000000000000000000000003008480010000000000000000000000000000000000000003008480010000000000000000000000000000000000000003008e80010000000000000000000000000015240000000003008e80010000000000000000000000000023240000010001009c05010000000000020000000000000000000000000003008e8001000000000000000000000000000000000000000300a48001000000000000000000000000000000000000000300a48001000000000000000000000000000000000000000300a68001000000000000000000000000000000000000000300aa8001000000000000000000000000000000000000000300aa8001000000000000000000000000000000000000000300b88001000000000000000000000000000000000000000300b88001000000000000000000000000000000000000000300b88001000000000000000000000000004f2400000000040048bc0100000000000000000000000000592400000000040050bc0100000000000000000000000000632400000000040058bc01000000000000000000000000006d24000002000300b880010000000000bc010000000000000000000000000300b88001000000000000000000000000000000000000000300b88001000000000000000000000000000000000000000300b88001000000000000000000000000000000000000000300ba8001000000000000000000000000000000000000000300d4800100000000000000000000000000d524000000000300de800100000000000000000000000000e324000000000300e6800100000000000000000000000000f124000000000300ee8001000000000000000000000000000000000000000300fe8001000000000000000000000000000000000000000300fe800100000000000000000000000000ff240000000003000681010000000000000000000000000000000000000003001681010000000000000000000000000000000000000003001681010000000000000000000000000000000000000003001a81010000000000000000000000000000000000000003001a81010000000000000000000000000000000000000003002481010000000000000000000000000000000000000003002481010000000000000000000000000000000000000003002881010000000000000000000000000000000000000003003681010000000000000000000000000000000000000003003681010000000000000000000000000000000000000003003e81010000000000000000000000000000000000000003003e81010000000000000000000000000000000000000003004881010000000000000000000000000000000000000003004881010000000000000000000000000000000000000003005081010000000000000000000000000000000000000003005081010000000000000000000000000000000000000003005681010000000000000000000000000000000000000003005681010000000000000000000000000000000000000003005a81010000000000000000000000000000000000000003005c81010000000000000000000000000000000000000003006881010000000000000000000000000000000000000003006a81010000000000000000000000000000000000000003007081010000000000000000000000000000000000000003007081010000000000000000000000000000000000000003007881010000000000000000000000000000000000000003007c81010000000000000000000000000000000000000003007c81010000000000000000000000000000000000000003008a81010000000000000000000000000000000000000003009081010000000000000000000000000000000000000003009481010000000000000000000000000000000000000003009481010000000000000000000000000000000000000003009881010000000000000000000000000000000000000003009881010000000000000000000000000000000000000003009e8101000000000000000000000000000000000000000300a08101000000000000000000000000000000000000000300a08101000000000000000000000000000000000000000300a28101000000000000000000000000000000000000000300a28101000000000000000000000000000000000000000300aa8101000000000000000000000000000000000000000300aa8101000000000000000000000000000000000000000300b48101000000000000000000000000000000000000000300b68101000000000000000000000000000000000000000300b68101000000000000000000000000000000000000000300b88101000000000000000000000000000000000000000300b88101000000000000000000000000000000000000000300c08101000000000000000000000000000000000000000300c08101000000000000000000000000000000000000000300c28101000000000000000000000000000000000000000300c88101000000000000000000000000000000000000000300c88101000000000000000000000000000000000000000300d48101000000000000000000000000000000000000000300d68101000000000000000000000000000000000000000300da8101000000000000000000000000000000000000000300da8101000000000000000000000000000000000000000300de8101000000000000000000000000000000000000000300e28101000000000000000000000000000000000000000300e88101000000000000000000000000000000000000000300e88101000000000000000000000000000000000000000300f48101000000000000000000000000000000000000000300fc8101000000000000000000000000000000000000000300fc8101000000000000000000000000000000000000000300fe81010000000000000000000000000000000000000003000082010000000000000000000000000000000000000003000882010000000000000000000000000000000000000003000882010000000000000000000000000000000000000003000a82010000000000000000000000000000000000000003000a82010000000000000000000000000000000000000003000e82010000000000000000000000000000000000000003000e82010000000000000000000000000000000000000003001282010000000000000000000000000000000000000003001282010000000000000000000000000000000000000003002682010000000000000000000000000000000000000003002c82010000000000000000000000000000000000000003003a8201000000000000000000000000000000000000000300428201000000000000000000000000000000000000000300428201000000000000000000000000000000000000000300468201000000000000000000000000000000000000000300468201000000000000000000000000000000000000000300568201000000000000000000000000000000000000000300708201000000000000000000000000000000000000000300748201000000000000000000000000000000000000000300748201000000000000000000000000000d250000020003007482010000000000b40000000000000000000000000003007482010000000000000000000000000000000000000003007482010000000000000000000000000000000000000003007482010000000000000000000000000000000000000003007682010000000000000000000000000000000000000003007882010000000000000000000000000000000000000003008082010000000000000000000000000000000000000003008282010000000000000000000000000000000000000003008282010000000000000000000000000000000000000003008682010000000000000000000000000000000000000003008682010000000000000000000000000000000000000003008e82010000000000000000000000000000000000000003008e8201000000000000000000000000000000000000000300948201000000000000000000000000000000000000000300948201000000000000000000000000000000000000000300988201000000000000000000000000000000000000000300a08201000000000000000000000000000000000000000300a48201000000000000000000000000000000000000000300b08201000000000000000000000000000000000000000300b08201000000000000000000000000000000000000000300b68201000000000000000000000000000000000000000300b68201000000000000000000000000000000000000000300ba8201000000000000000000000000000000000000000300c28201000000000000000000000000000000000000000300c88201000000000000000000000000000000000000000300d08201000000000000000000000000000000000000000300d48201000000000000000000000000000000000000000300e08201000000000000000000000000000000000000000300e68201000000000000000000000000000000000000000300ee8201000000000000000000000000000000000000000300f48201000000000000000000000000000000000000000300fc82010000000000000000000000000000000000000003000283010000000000000000000000000000000000000003000a83010000000000000000000000000000000000000003000e83010000000000000000000000000000000000000003001883010000000000000000000000000000000000000003001883010000000000000000000000000000000000000003002283010000000000000000000000000000000000000003002483010000000000000000000000000000000000000003002883010000000000000000000000000000000000000003002883010000000000000000000000000040250000020003002883010000000000380000000000000000000000000003002883010000000000000000000000000000000000000003002883010000000000000000000000000000000000000003002883010000000000000000000000000000000000000003002a83010000000000000000000000000000000000000003002a83010000000000000000000000000000000000000003002c8301000000000000000000000000007125000000000300468301000000000000000000000000007f250000010001006806010000000000300000000000000000000000000003005a83010000000000000000000000000000000000000003005c830100000000000000000000000000000000000000030060830100000000000000000000000000000000000000030060830100000000000000000000000000ab2500000200030060830100000000000a0000000000000000000000000003006083010000000000000000000000000000000000000003006083010000000000000000000000000000000000000003006083010000000000000000000000000000000000000003006083010000000000000000000000000000000000000003006a83010000000000000000000000000000000000000003006a83010000000000000000000000000001260000020003006a83010000000000b60000000000000000000000000003006a83010000000000000000000000000000000000000003006a83010000000000000000000000000000000000000003006a83010000000000000000000000000000000000000003006c83010000000000000000000000000000000000000003006c83010000000000000000000000000000000000000003006e83010000000000000000000000000000000000000003007883010000000000000000000000000000000000000003007883010000000000000000000000000000000000000003007a83010000000000000000000000000000000000000003007a83010000000000000000000000000000000000000003007e83010000000000000000000000000000000000000003007e83010000000000000000000000000000000000000003008683010000000000000000000000000000000000000003008683010000000000000000000000000000000000000003008c83010000000000000000000000000000000000000003008c83010000000000000000000000000000000000000003009083010000000000000000000000000000000000000003009883010000000000000000000000000000000000000003009c8301000000000000000000000000000000000000000300a88301000000000000000000000000000000000000000300a88301000000000000000000000000000000000000000300ae8301000000000000000000000000000000000000000300ae8301000000000000000000000000000000000000000300b28301000000000000000000000000000000000000000300ba8301000000000000000000000000000000000000000300c08301000000000000000000000000000000000000000300c88301000000000000000000000000000000000000000300cc8301000000000000000000000000000000000000000300d88301000000000000000000000000000000000000000300de8301000000000000000000000000000000000000000300e68301000000000000000000000000000000000000000300ec8301000000000000000000000000000000000000000300f48301000000000000000000000000000000000000000300fa83010000000000000000000000000000000000000003000284010000000000000000000000000000000000000003000684010000000000000000000000000000000000000003001084010000000000000000000000000000000000000003001084010000000000000000000000000000000000000003001a84010000000000000000000000000000000000000003001a84010000000000000000000000000000000000000003001c840100000000000000000000000000000000000000030020840100000000000000000000000000000000000000030020840100000000000000000000000000592600000200030020840100000000003a00000000000000000000000000030020840100000000000000000000000000000000000000030020840100000000000000000000000000000000000000030020840100000000000000000000000000000000000000030022840100000000000000000000000000000000000000030022840100000000000000000000000000000000000000030024840100000000000000000000000000af260000000003004084010000000000000000000000000000000000000003004084010000000000000000000000000000000000000003004084010000000000000000000000000000000000000003005484010000000000000000000000000000000000000003005484010000000000000000000000000000000000000003005684010000000000000000000000000000000000000003005a84010000000000000000000000000000000000000003005a840100000000000000000000000000bd260000020003005a84010000000000200100000000000000000000000003005a84010000000000000000000000000000000000000003005a84010000000000000000000000000000000000000003005a84010000000000000000000000000000000000000003005c84010000000000000000000000000000000000000003006a84010000000000000000000000000000000000000003006c84010000000000000000000000000000000000000003007084010000000000000000000000000000000000000003007084010000000000000000000000000000000000000003007284010000000000000000000000000000000000000003007284010000000000000000000000000000000000000003007a84010000000000000000000000000000000000000003007e84010000000000000000000000000000000000000003007e84010000000000000000000000000000000000000003008284010000000000000000000000000000000000000003008284010000000000000000000000000000000000000003008684010000000000000000000000000000000000000003008684010000000000000000000000000000000000000003008a84010000000000000000000000000000000000000003008a84010000000000000000000000000000000000000003008e84010000000000000000000000000000000000000003008e840100000000000000000000000000000000000000030090840100000000000000000000000000000000000000030094840100000000000000000000000000f926000000000300988401000000000000000000000000000727000001000100960501000000000002000000000000000000000000000300988401000000000000000000000000000000000000000300a28401000000000000000000000000000000000000000300a68401000000000000000000000000000000000000000300a68401000000000000000000000000003327000000000300b08401000000000000000000000000004127000001000100980501000000000002000000000000000000000000000300bc8401000000000000000000000000000000000000000300bc8401000000000000000000000000000000000000000300be8401000000000000000000000000006d27000000000300c48401000000000000000000000000007b270000010001009a0501000000000001000000000000000000000000000300cc8401000000000000000000000000000000000000000300cc8401000000000000000000000000000000000000000300d68401000000000000000000000000000000000000000300d68401000000000000000000000000000000000000000300d88401000000000000000000000000000000000000000300d88401000000000000000000000000000000000000000300dc8401000000000000000000000000000000000000000300dc8401000000000000000000000000000000000000000300de8401000000000000000000000000000000000000000300de8401000000000000000000000000000000000000000300ea8401000000000000000000000000000000000000000300ea8401000000000000000000000000000000000000000300ee8401000000000000000000000000000000000000000300ee8401000000000000000000000000000000000000000300f08401000000000000000000000000000000000000000300f48401000000000000000000000000000000000000000300f48401000000000000000000000000000000000000000300fc8401000000000000000000000000000000000000000300fc84010000000000000000000000000000000000000003000685010000000000000000000000000000000000000003000685010000000000000000000000000000000000000003000a85010000000000000000000000000000000000000003000e85010000000000000000000000000000000000000003001685010000000000000000000000000000000000000003001e850100000000000000000000000000000000000000030032850100000000000000000000000000000000000000030032850100000000000000000000000000000000000000030036850100000000000000000000000000a72700000000030036850100000000000000000000000000b52700000100010058050100000000003000000000000000000000000000030036850100000000000000000000000000000000000000030040850100000000000000000000000000000000000000030040850100000000000000000000000000000000000000030048850100000000000000000000000000000000000000030048850100000000000000000000000000e1270000000003004e850100000000000000000000000000ef270000010001009405010000000000020000000000000000000000000003005a85010000000000000000000000000000000000000003005a85010000000000000000000000000000000000000003005c85010000000000000000000000000000000000000003005c85010000000000000000000000000000000000000003006085010000000000000000000000000000000000000003006685010000000000000000000000000000000000000003007685010000000000000000000000000000000000000003007a85010000000000000000000000000000000000000003007a85010000000000000000000000000000000000000003007a85010000000000000000000000000000000000000003007a85010000000000000000000000000000000000000003007a85010000000000000000000000000000000000000003007c85010000000000000000000000000000000000000003008485010000000000000000000000000000000000000003008685010000000000000000000000000000000000000003008685010000000000000000000000000000000000000003009285010000000000000000000000000000000000000003009285010000000000000000000000000000000000000003009e85010000000000000000000000000000000000000003009e8501000000000000000000000000000000000000000300ac8501000000000000000000000000000000000000000300ac8501000000000000000000000000000000000000000300ae8501000000000000000000000000000000000000000300b28501000000000000000000000000000000000000000300b48501000000000000000000000000000000000000000300b68501000000000000000000000000000000000000000300b68501000000000000000000000000000000000000000300b88501000000000000000000000000000000000000000300b88501000000000000000000000000000000000000000300c28501000000000000000000000000000000000000000300c48501000000000000000000000000000000000000000300cc8501000000000000000000000000000000000000000300cc8501000000000000000000000000000000000000000300d28501000000000000000000000000000000000000000300d28501000000000000000000000000000000000000000300d48501000000000000000000000000000000000000000300d48501000000000000000000000000001b28000000000300da85010000000000000000000000000029280000010001009b0501000000000001000000000000000000000000000300e88501000000000000000000000000000000000000000300e88501000000000000000000000000000000000000000300ea8501000000000000000000000000000000000000000300ea8501000000000000000000000000005528000000000300f085010000000000000000000000000063280000010001003a05010000000000010000000000000000000000000003000086010000000000000000000000000000000000000003000086010000000000000000000000000000000000000003000486010000000000000000000000000000000000000003000486010000000000000000000000000000000000000003000e8601000000000000000000000000000000000000000300128601000000000000000000000000000000000000000300128601000000000000000000000000000000000000000300128601000000000000000000000000000000000000000300128601000000000000000000000000000000000000000300128601000000000000000000000000000000000000000300148601000000000000000000000000000000000000000300148601000000000000000000000000000000000000000300168601000000000000000000000000000000000000000300208601000000000000000000000000000000000000000300208601000000000000000000000000008f2800000200030020860100000000001600000000000000000000000000030020860100000000000000000000000000000000000000030020860100000000000000000000000000d72800000000030020860100000000000000000000000000000000000000030020860100000000000000000000000000e5280000010001009806010000000000020000000000000000000000000003002086010000000000000000000000000000000000000003003686010000000000000000000000000000000000000003003686010000000000000000000000000000000000000003003686010000000000000000000000000011290000020003003686010000000000a20000000000000000000000000003003686010000000000000000000000000000000000000003003686010000000000000000000000000000000000000003003686010000000000000000000000000000000000000003003886010000000000000000000000000000000000000003003e8601000000000000000000000000000000000000000300408601000000000000000000000000000000000000000300408601000000000000000000000000000000000000000300428601000000000000000000000000000000000000000300428601000000000000000000000000000000000000000300448601000000000000000000000000000000000000000300448601000000000000000000000000007229000000000300488601000000000000000000000000008029000001000100c0060100000000001100000000000000000000000000030054860100000000000000000000000000000000000000030054860100000000000000000000000000000000000000030060860100000000000000000000000000ac2900000000030060860100000000000000000000000000ba29000001000100a006010000000000200000000000000000000000000003006086010000000000000000000000000000000000000003007486010000000000000000000000000000000000000003007486010000000000000000000000000000000000000003007686010000000000000000000000000000000000000003007a86010000000000000000000000000000000000000003007c86010000000000000000000000000000000000000003007e86010000000000000000000000000000000000000003007e86010000000000000000000000000000000000000003008086010000000000000000000000000000000000000003008086010000000000000000000000000000000000000003008a86010000000000000000000000000000000000000003008c86010000000000000000000000000000000000000003009486010000000000000000000000000000000000000003009486010000000000000000000000000000000000000003009a86010000000000000000000000000000000000000003009a86010000000000000000000000000000000000000003009c86010000000000000000000000000000000000000003009c860100000000000000000000000000e629000000000300a28601000000000000000000000000000000000000000300b08601000000000000000000000000000000000000000300b08601000000000000000000000000000000000000000300b28601000000000000000000000000000000000000000300b2860100000000000000000000000000f429000000000300b88601000000000000000000000000000000000000000300c88601000000000000000000000000000000000000000300c88601000000000000000000000000000000000000000300cc8601000000000000000000000000000000000000000300cc8601000000000000000000000000000000000000000300d48601000000000000000000000000000000000000000300d88601000000000000000000000000000000000000000300d8860100000000000000000000000000022a000002000300d88601000000000070000000000000000000000000000300d88601000000000000000000000000000000000000000300d88601000000000000000000000000000000000000000300d88601000000000000000000000000000000000000000300da8601000000000000000000000000000000000000000300dc8601000000000000000000000000000000000000000300de8601000000000000000000000000000000000000000300de8601000000000000000000000000000000000000000300e68601000000000000000000000000000000000000000300e68601000000000000000000000000000000000000000300ee8601000000000000000000000000000000000000000300ee8601000000000000000000000000000000000000000300f08601000000000000000000000000000000000000000300f08601000000000000000000000000000000000000000300f48601000000000000000000000000000000000000000300f48601000000000000000000000000000000000000000300fc8601000000000000000000000000000000000000000300fe8601000000000000000000000000000000000000000300fe86010000000000000000000000000000000000000003000687010000000000000000000000000000000000000003000687010000000000000000000000000000000000000003000a87010000000000000000000000000000000000000003000a87010000000000000000000000000000000000000003001487010000000000000000000000000000000000000003001487010000000000000000000000000000000000000003001e870100000000000000000000000000622a0000000003001e87010000000000000000000000000000000000000003001e87010000000000000000000000000000000000000003003487010000000000000000000000000000000000000003003487010000000000000000000000000000000000000003003687010000000000000000000000000000000000000003003a87010000000000000000000000000000000000000003003a870100000000000000000000000000000000000000030048870100000000000000000000000000000000000000030048870100000000000000000000000000000000000000030048870100000000000000000000000000702a0000020003004887010000000000520000000000000000000000000003004887010000000000000000000000000000000000000003004a8701000000000000000000000000000000000000000300548701000000000000000000000000001c2b0000020003009a870100000000007e0000000000000000000000000003009a87010000000000000000000000000000000000000003009a87010000000000000000000000000000000000000003009c8701000000000000000000000000000000000000000300a287010000000000000000000000000000000000000003001888010000000000000000000000000000000000000003001888010000000000000000000000000000000000000003001a880100000000000000000000000000000000000000030022880100000000000000000000000000762b000002000300b691010000000000080000000000000000000000000003007a880100000000000000000000000000852b0000020003007a88010000000000300000000000000000000000000003007a8801000000000000000000000000000000000000000300aa8801000000000000000000000000000000000000000300aa8801000000000000000000000000000000000000000300ac8801000000000000000000000000000000000000000300b0880100000000000000000000000000cd2b000002000300be9101000000000008000000000000000000000000000300f8880100000000000000000000000000e12b000002000300f88801000000000068000000000000000000000000000300f88801000000000000000000000000000000000000000300fa880100000000000000000000000000000000000000030004890100000000000000000000000000222c00000200030060890100000000007e000000000000000000000000000300608901000000000000000000000000000000000000000300608901000000000000000000000000000000000000000300628901000000000000000000000000000000000000000300688901000000000000000000000000007c2c000002000300de8901000000000052000000000000000000000000000300de8901000000000000000000000000000000000000000300de8901000000000000000000000000000000000000000300e08901000000000000000000000000000000000000000300e68901000000000000000000000000000000000000000300308a01000000000000000000000000000000000000000300308a01000000000000000000000000000000000000000300328a01000000000000000000000000000000000000000300368a01000000000000000000000000000000000000000300868a0100000000000000000000000000af2c000002000300868a01000000000082010000000000000000000000000300868a01000000000000000000000000000000000000000300888a01000000000000000000000000000000000000000300968a0100000000000000000000000000e02c000000000300688b0100000000000000000000000000ee2c000001000100a0070100000000001c00000000000000f82c000000000300728b0100000000000000000000000000062d0000000003007c8b0100000000000000000000000000142d000000000300908b0100000000000000000000000000222d000000000300988b0100000000000000000000000000302d000001000100f80601000000000020000000000000005a2d000000000300a68b0100000000000000000000000000682d00000100010006080100000000002f00000000000000932d000000000300b48b0100000000000000000000000000a12d00000100010035080100000000003200000000000000cc2d000000000300ce8b0100000000000000000000000000da2d000000000300d68b0100000000000000000000000000e82d00000100010080070100000000002000000000000000122e000000000300f08b0100000000000000000000000000202e000001000100bc070100000000001c000000000000004b2e000000000300fa8b0100000000000000000000000000592e000001000100d8070100000000002e000000000000000000000000000300088c0100000000000000000000000000842e000002000300088c01000000000028000000000000000000000000000300088c0100000000000000000000000000df2e0000000003000e8c0100000000000000000000000000ed2e000001000100280a0100000000005000000000000000572f000000000300188c0100000000000000000000000000652f000001000100780a01000000000050000000000000000000000000000300308c0100000000000000000000000000d32f000002000300308c01000000000062000000000000000000000000000300308c01000000000000000000000000000000000000000300328c01000000000000000000000000000c30000000000300528c01000000000000000000000000001a300000000003005e8c01000000000000000000000000002830000001000100180701000000000018000000000000005230000000000300668c01000000000000000000000000006030000001000100300701000000000020000000000000008a300000000003007c8c01000000000000000000000000009830000001000100670801000000000026000000000000000000000000000300928c0100000000000000000000000000c330000002000300928c01000000000068000000000000000000000000000300928c01000000000000000000000000000000000000000300948c01000000000000000000000000000000000000000300988c01000000000000000000000000000231000000000300c48c01000000000000000000000000001031000000000300cc8c01000000000000000000000000001e31000000000300e68c01000000000000000000000000002c310000010001008d080100000000000d000000000000000000000000000300fa8c01000000000000000000000000000000000000000300fa8c01000000000000000000000000000000000000000300fc8c01000000000000000000000000000000000000000300008d01000000000000000000000000005731000000000300388d010000000000000000000000000000000000000003004e8d010000000000000000000000000000000000000003004e8d01000000000000000000000000000000000000000300508d01000000000000000000000000000000000000000300628d01000000000000000000000000006531000000000300e88d01000000000000000000000000007331000000000300768e01000000000000000000000000008131000000000300808e01000000000000000000000000008f310000010001009a080100000000000e00000000000000ba310000000003008c8e0100000000000000000000000000c831000000000300968e0100000000000000000000000000d631000000000300a08e0100000000000000000000000000e431000000000300aa8e0100000000000000000000000000f231000000000300b48e01000000000000000000000000000000000000000300ca8e01000000000000000000000000000000000000000300ca8e01000000000000000000000000000000000000000300cc8e01000000000000000000000000000000000000000300d28e010000000000000000000000000000320000000003000c8f01000000000000000000000000000e32000000000300148f01000000000000000000000000001c320000000003002e8f01000000000000000000000000002a32000001000100a8080100000000000e000000000000000000000000000300428f01000000000000000000000000000000000000000300428f01000000000000000000000000000000000000000300448f010000000000000000000000000000000000000003004a8f010000000000000000000000000055320000000003008a8f01000000000000000000000000006332000000000300928f01000000000000000000000000007132000000000300ac8f01000000000000000000000000007f32000001000100b6080100000000000d000000000000000000000000000300c08f01000000000000000000000000000000000000000300c08f01000000000000000000000000000000000000000300c28f01000000000000000000000000000000000000000300ca8f0100000000000000000000000000aa320000000003002c900100000000000000000000000000b83200000000030034900100000000000000000000000000c6320000000003004e900100000000000000000000000000d432000001000100c3080100000000001200000000000000000000000000030062900100000000000000000000000000ff3200000200030062900100000000007a0000000000000000000000000003006290010000000000000000000000000000000000000003006490010000000000000000000000000000000000000003006a9001000000000000000000000000006333000000000300ba9001000000000000000000000000000000000000000300dc9001000000000000000000000000000000000000000300dc9001000000000000000000000000000000000000000300de9001000000000000000000000000000000000000000300ea9001000000000000000000000000007133000000000300449101000000000000000000000000007f33000001000100d8080100000000002000000000000000000000000000030096910100000000000000000000000000aa33000002000300969101000000000010000000000000000000000000000300969101000000000000000000000000000000000000000300a69101000000000000000000000000000000000000000300a69101000000000000000000000000000000000000000300ae9101000000000000000000000000000000000000000300ae9101000000000000000000000000000000000000000300b69101000000000000000000000000000000000000000300b69101000000000000000000000000000000000000000300be9101000000000000000000000000000000000000000300be9101000000000000000000000000000000000000000300c69101000000000000000000000000000000000000000300c69101000000000000000000000000000000000000000300d09101000000000000000000000000000000000000000300d09101000000000000000000000000000000000000000300d29101000000000000000000000000000000000000000300da910100000000000000000000000000fb330000000003002492010000000000000000000000000000000000000003004292010000000000000000000000000009340000020003004292010000000000ca020000000000000000000000000300429201000000000000000000000000000000000000000300449201000000000000000000000000000000000000000300549201000000000000000000000000009334000000000300ce940100000000000000000000000000a134000000000300e2940100000000000000000000000000af34000000000300ec940100000000000000000000000000bd34000000000300f494010000000000000000000000000000000000000003000c95010000000000000000000000000000000000000003000c950100000000000000000000000000cb340000000003000e950100000000000000000000000000d93400000000010088010100000000000000000000000000e4340000000003001e950100000000000000000000000000ee3400000000030020950100000000000000000000000000f834000000000300229501000000000000000000000000000235000000000300269501000000000000000000000000000c350000000003002a95010000000000000000000000000000000000000003003495010000000000000000000000000000000000000003003495010000000000000000000000000000000000000003003695010000000000000000000000000000000000000003004695010000000000000000000000000000000000000003009896010000000000000000000000000000000000000003009896010000000000000000000000000000000000000003009c9601000000000000000000000000000000000000000300c09601000000000000000000000000001635000000000300209a01000000000000000000000000002435000000000300a29b0100000000000000000000000000323500000100010030040100000000001c000000000000003b35000000000300ac9b01000000000000000000000000004935000000000300b69b01000000000000000000000000005735000000000300c09b01000000000000000000000000006535000000000300ca9b01000000000000000000000000007335000000000300de9b01000000000000000000000000008135000000000300e69b01000000000000000000000000008f350000010001009009010000000000200000000000000000000000000003001e9c010000000000000000000000000000000000000003001e9c01000000000000000000000000000000000000000300209c01000000000000000000000000000000000000000300369c0100000000000000000000000000ba35000000000300f49e0100000000000000000000000000c835000000000300089f0100000000000000000000000000d635000001000100d0090100000000002b000000000000000236000000000300169f010000000000000000000000000010360000000003001e9f01000000000000000000000000000000000000000300369f01000000000000000000000000000000000000000300369f01000000000000000000000000000000000000000300389f010000000000000000000000000000000000000003003e9f01000000000000000000000000000000000000000300c89f01000000000000000000000000000000000000000300c89f01000000000000000000000000000000000000000300ca9f01000000000000000000000000000000000000000300e49f01000000000000000000000000001e360000000003001ca301000000000000000000000000002c3600000000030030a301000000000000000000000000003a3600000000030038a30100000000000000000000000000483600000000030050a301000000000000000000000000005636000001000100fb090100000000002900000000000000000000000000030068a30100000000000000000000000000000000000000030068a3010000000000000000000000000000000000000003006aa30100000000000000000000000000000000000000030076a301000000000000000000000000008236000000000300c8a401000000000000000000000000000000000000000300eea40100000000000000000000000000903600000100060018bd0100000000000010080000000000bb3600000100060018cd0900000000000010000000000000ec360000010001007c0301000000000023000000000000001737000001000100b00301000000000033000000000000004237000001000100f8080100000000000a000000000000006d3700000100010002090100000000000a0000000000000098370000010001000c090100000000000b00000000000000c33700000100010017090100000000000600000000000000ee370000010001001d09010000000000060000000000000019380000010001002309010000000000090000000000000044380000010001002c0901000000000006000000000000000000000000000800000000000000000000000000000000000000000000000b006f2900000000000000000000000000000000000000000b00114300000000000000000000000000006f38000000000f00000000000000000000000000000000000000000000000b00051200000000000000000000000000000000000000000a00700e00000000000000000000000000000000000000000b001e2d00000000000000000000000000000000000000000b00000000000000000000000000000000000000000000000b00c44b00000000000000000000000000000000000000000b00783500000000000000000000000000000000000000000b00463c00000000000000000000000000000000000000000b001d0e00000000000000000000000000000000000000000800740000000000000000000000000000000000000000000b00f91500000000000000000000000000008338000000000f00880000000000000000000000000000000000000000000a00a00e00000000000000000000000000000000000000000b00da1800000000000000000000000000000000000000000b001f0500000000000000000000000000000000000000000b007d0c00000000000000000000000000000000000000000b002f1600000000000000000000000000000000000000000b00f03200000000000000000000000000000000000000000b002b0c00000000000000000000000000000000000000000b005c3c00000000000000000000000000000000000000000b00ab3000000000000000000000000000000000000000000b00fa3500000000000000000000000000000000000000000b00712300000000000000000000000000000000000000000b00942800000000000000000000000000000000000000000b00c52100000000000000000000000000000000000000000b00e52a00000000000000000000000000000000000000000b00194600000000000000000000000000000000000000000b006b3800000000000000000000000000000000000000000b00833700000000000000000000000000000000000000000b00c50b00000000000000000000000000000000000000000b00f90300000000000000000000000000000000000000000b00ad0c00000000000000000000000000000000000000000b005f3f00000000000000000000000000000000000000000b00c43000000000000000000000000000000000000000000b002c1700000000000000000000000000000000000000000b004d0b00000000000000000000000000000000000000000b00e93400000000000000000000000000000000000000000b00a60000000000000000000000000000000000000000000b00c14600000000000000000000000000000000000000000b00d71200000000000000000000000000000000000000000b00084100000000000000000000000000000000000000000b006c4500000000000000000000000000000000000000000b002b0500000000000000000000000000000000000000000b00060800000000000000000000000000000000000000000b00cc0000000000000000000000000000000000000000000b00052800000000000000000000000000000000000000000b00a73000000000000000000000000000000000000000000b00351200000000000000000000000000000000000000000b00a43100000000000000000000000000000000000000000b00454800000000000000000000000000000000000000000b004e2700000000000000000000000000000000000000000b002c3e00000000000000000000000000000000000000000b00101300000000000000000000000000000000000000000b00104600000000000000000000000000000000000000000b00403b00000000000000000000000000000000000000000b009c4800000000000000000000000000000000000000000b00632e00000000000000000000000000000000000000000b009b1500000000000000000000000000000000000000000b008a3500000000000000000000000000000000000000000a00000000000000000000000000000000000000000000000a00400000000000000000000000000000000000000000000a00700000000000000000000000000000000000000000000a00a00000000000000000000000000000000000000000000b00a30b00000000000000000000000000000000000000000b00412b00000000000000000000000000000000000000000b00713b00000000000000000000000000000000000000000b00be2d00000000000000000000000000000000000000000b00482900000000000000000000000000000000000000000b00242900000000000000000000000000000000000000000b00db1300000000000000000000000000000000000000000b00b11b00000000000000000000000000000000000000000b003c4400000000000000000000000000000000000000000b000d4700000000000000000000000000000000000000000b00ce3800000000000000000000000000000000000000000b00501400000000000000000000000000000000000000000b00032e00000000000000000000000000000000000000000a00200900000000000000000000000000000000000000000a00500900000000000000000000000000000000000000000a00800900000000000000000000000000000000000000000a00b00900000000000000000000000000000000000000000a00e00900000000000000000000000000000000000000000b00650700000000000000000000000000000000000000000b00873200000000000000000000000000000000000000000b006f0700000000000000000000000000000000000000000b001f0300000000000000000000000000000000000000000a00800d00000000000000000000000000000000000000000a00b00d00000000000000000000000000000000000000000a00e00d00000000000000000000000000000000000000000a00100e00000000000000000000000000000000000000000a00400e00000000000000000000000000000000000000000b001f4a00000000000000000000000000000000000000000b00370a00000000000000000000000000000000000000000b006c0a00000000000000000000000000000000000000000b007f0300000000000000000000000000000000000000000b00672e00000000000000000000000000000000000000000b00114900000000000000000000000000000000000000000b00f44000000000000000000000000000000000000000000b00b90c00000000000000000000000000000000000000000b00230500000000000000000000000000000000000000000b00890200000000000000000000000000000000000000000b00e03100000000000000000000000000000000000000000a00d00000000000000000000000000000000000000000000a00100100000000000000000000000000000000000000000a00400100000000000000000000000000000000000000000a00700100000000000000000000000000000000000000000a00a00100000000000000000000000000000000000000000a00d00100000000000000000000000000000000000000000a00000200000000000000000000000000000000000000000a00300200000000000000000000000000000000000000000a00800200000000000000000000000000000000000000000b00c04700000000000000000000000000000000000000000b00f92d00000000000000000000000000000000000000000a00b00200000000000000000000000000000000000000000a00e00200000000000000000000000000000000000000000a00100300000000000000000000000000000000000000000a00400300000000000000000000000000000000000000000a00700300000000000000000000000000000000000000000a00a00300000000000000000000000000000000000000000a00d00300000000000000000000000000000000000000000a00000400000000000000000000000000000000000000000a00300400000000000000000000000000000000000000000a00800400000000000000000000000000000000000000000a00b00400000000000000000000000000000000000000000a00000500000000000000000000000000000000000000000a00300500000000000000000000000000000000000000000a00800500000000000000000000000000000000000000000a00b00500000000000000000000000000000000000000000a00f00500000000000000000000000000000000000000000a00600600000000000000000000000000000000000000000a00b00600000000000000000000000000000000000000000a00f00600000000000000000000000000000000000000000a00200700000000000000000000000000000000000000000a00500700000000000000000000000000000000000000000b003c3800000000000000000000000000000000000000000b00ae2d00000000000000000000000000000000000000000b00371700000000000000000000000000000000000000000b00372b00000000000000000000000000000000000000000b00263100000000000000000000000000000000000000000b00172900000000000000000000000000000000000000000b001a2700000000000000000000000000000000000000000b00431c00000000000000000000000000000000000000000b001f0700000000000000000000000000000000000000000b00572300000000000000000000000000000000000000000b001e1a00000000000000000000000000000000000000000b00f81600000000000000000000000000000000000000000b00fb2e00000000000000000000000000000000000000000b00012f00000000000000000000000000000000000000000b00cf4900000000000000000000000000000000000000000b00d81900000000000000000000000000000000000000000b00fa0800000000000000000000000000000000000000000b008b4900000000000000000000000000000000000000000b001b0f00000000000000000000000000000000000000000b001f0900000000000000000000000000000000000000000b00453900000000000000000000000000000000000000000a00800700000000000000000000000000000000000000000a00b00700000000000000000000000000000000000000000a00e00700000000000000000000000000000000000000000a00100800000000000000000000000000000000000000000a00400800000000000000000000000000000000000000000a00700800000000000000000000000000000000000000000a00a00800000000000000000000000000000000000000000a00e00800000000000000000000000000000000000000000b00f10100000000000000000000000000000000000000000b00d53c00000000000000000000000000000000000000000b00bd3800000000000000000000000000000000000000000b00ec3700000000000000000000000000000000000000000b00923500000000000000000000000000000000000000000a00100a00000000000000000000000000000000000000000a00400a00000000000000000000000000000000000000000a00700a00000000000000000000000000000000000000000a00a00a00000000000000000000000000000000000000000a00d00a00000000000000000000000000000000000000000a00000b00000000000000000000000000000000000000000b00623d00000000000000000000000000000000000000000b00f64400000000000000000000000000000000000000000b00920400000000000000000000000000000000000000000b00d11900000000000000000000000000000000000000000b00fc2200000000000000000000000000000000000000000b003d2900000000000000000000000000000000000000000b008f4900000000000000000000000000000000000000000b00ae4600000000000000000000000000000000000000000b00bd0900000000000000000000000000000000000000000a00b00b00000000000000000000000000000000000000000a00e00b00000000000000000000000000000000000000000a00100c00000000000000000000000000000000000000000a00400c00000000000000000000000000000000000000000a00700c00000000000000000000000000000000000000000a00b00c00000000000000000000000000000000000000000b00bd1c00000000000000000000000000000000000000000b00b54700000000000000000000000000000000000000000b00821c00000000000000000000000000000000000000000b00b92d00000000000000000000000000000000000000000b00f10800000000000000000000000000000000000000000b001f3500000000000000000000000000000000000000000b00693100000000000000000000000000000000000000000b00ec2200000000000000000000000000000000000000000b00e82f00000000000000000000000000000000000000000a00300b00000000000000000000000000000000000000000b004d1800000000000000000000000000000000000000000b00ee2f00000000000000000000000000000000000000000b00c54400000000000000000000000000000000000000000b00994b00000000000000000000000000000000000000000b00ef4700000000000000000000000000000000000000000b00284200000000000000000000000000000000000000000b00534200000000000000000000000000000000000000000a00700b00000000000000000000000000000000000000000b00963700000000000000000000000000000000000000000b00780900000000000000000000000000000000000000000b00b40f00000000000000000000000000000000000000000b00210c00000000000000000000000000000000000000000b005f3000000000000000000000000000000000000000000b00ff0f00000000000000000000000000000000000000000b008c3900000000000000000000000000000000000000000b00164a00000000000000000000000000000000000000000b00954800000000000000000000000000000000000000000b00820900000000000000000000000000000000000000000b00fd4b00000000000000000000000000000000000000000b00903900000000000000000000000000000000000000000b00f90900000000000000000000000000000000000000000b00681000000000000000000000000000000000000000000b00b13100000000000000000000000000000000000000000b00fa1c00000000000000000000000000000000000000000b00792300000000000000000000000000000000000000000b007a3300000000000000000000000000000000000000000b00564500000000000000000000000000000000000000000b00c63a00000000000000000000000000000000000000000b00c10100000000000000000000000000000000000000000b006b2a00000000000000000000000000000000000000000b00274100000000000000000000000000000000000000000b00b34a00000000000000000000000000000000000000000b000b3e00000000000000000000000000000000000000000b00f91a00000000000000000000000000000000000000000b00b73c00000000000000000000000000000000000000000b004c3600000000000000000000000000000000000000000b00120000000000000000000000000000000000000000000b00fd1900000000000000000000000000000000000000000b002b2d00000000000000000000000000000000000000000b00514900000000000000000000000000000000000000000b00f53100000000000000000000000000000000000000000b00d52100000000000000000000000000000000000000000b00e52100000000000000000000000000000000000000000b005f3400000000000000000000000000000000000000000b00a94a00000000000000000000000000000000000000000b00033700000000000000000000000000000000000000000b00c20a00000000000000000000000000000000000000000b00b03a00000000000000000000000000000000000000000b009b0b00000000000000000000000000000000000000000b00731b00000000000000000000000000000000000000000b00dd4100000000000000000000000000000000000000000b00641100000000000000000000000000000000000000000b002a1a00000000000000000000000000000000000000000b00a91a00000000000000000000000000000000000000000b00f62700000000000000000000000000000000000000000b00f14300000000000000000000000000000000000000000b00e24600000000000000000000000000000000000000000b00852500000000000000000000000000000000000000000b00ac3d00000000000000000000000000000000000000000b00b30500000000000000000000000000000000000000000b00c33d00000000000000000000000000000000000000000b00434100000000000000000000000000000000000000000b00b00800000000000000000000000000000000000000000b00342800000000000000000000000000000000000000000b00802800000000000000000000000000000000000000000b00f53700000000000000000000000000000000000000000b009f3a00000000000000000000000000000000000000000b00531900000000000000000000000000000000000000000b00ab1100000000000000000000000000000000000000000b00974100000000000000000000000000000000000000000b00432f00000000000000000000000000000000000000000b001f2600000000000000000000000000000000000000000b00280900000000000000000000000000000000000000000b00a90d00000000000000000000000000000000000000000b00ca1700000000000000000000000000000000000000000b004c0400000000000000000000000000000000000000000b00a91900000000000000000000000000000000000000000b000f0700000000000000000000000000000000000000000b00ab4200000000000000000000000000000000000000000b007a3900000000000000000000000000000000000000000b00b40300000000000000000000000000000000000000000b004a0500000000000000000000000000000000000000000b00ed3100000000000000000000000000000000000000000b00753400000000000000000000000000000000000000000b00f02800000000000000000000000000000000000000000b00400d00000000000000000000000000000000000000000b00d91100000000000000000000000000000000000000000b00353e00000000000000000000000000000000000000000b00123100000000000000000000000000000000000000000b008d3700000000000000000000000000000000000000000b00fa0100000000000000000000000000000000000000000b00364600000000000000000000000000000000000000000b00542f00000000000000000000000000000000000000000b006c1700000000000000000000000000000000000000000b00c31400000000000000000000000000000000000000000b00ec0c00000000000000000000000000000000000000000b00594900000000000000000000000000000000000000000b005a1400000000000000000000000000000000000000000b00983b00000000000000000000000000000000000000000b00b71b00000000000000000000000000000000000000000b00573d00000000000000000000000000000000000000000b00b22d00000000000000000000000000000000000000000b00d81700000000000000000000000000000000000000000b00a63b00000000000000000000000000000000000000000b00de3b00000000000000000000000000000000000000000b00744700000000000000000000000000000000000000000b00341c00000000000000000000000000000000000000000b00760f00000000000000000000000000000000000000000b00a93e00000000000000000000000000000000000000000b00242d00000000000000000000000000000000000000000b00b02900000000000000000000000000000000000000000b00494300000000000000000000000000000000000000000b00381200000000000000000000000000000000000000000b00842300000000000000000000000000000000000000000b00663c00000000000000000000000000000000000000000b00ad3f00000000000000000000000000000000000000000b008f3600000000000000000000000000000000000000000b00f60000000000000000000000000000000000000000000b003a0800000000000000000000000000000000000000000b00ba0e00000000000000000000000000000000000000000b00801000000000000000000000000000000000000000000b00861000000000000000000000000000000000000000000b005a2700000000000000000000000000000000000000000b009b3900000000000000000000000000000000000000000b00b50c00000000000000000000000000000000000000000b00804000000000000000000000000000000000000000000b00901000000000000000000000000000000000000000000b00b84600000000000000000000000000000000000000000b00712e00000000000000000000000000000000000000000b00752e00000000000000000000000000000000000000000b00ff1c00000000000000000000000000000000000000000b00304a00000000000000000000000000000000000000000b005e4300000000000000000000000000000000000000000b001c1f00000000000000000000000000000000000000000b00294a00000000000000000000000000000000000000000b00790700000000000000000000000000000000000000000b00781200000000000000000000000000000000000000000b000c0000000000000000000000000000000000000000000b005f4500000000000000000000000000000000000000000b00441600000000000000000000000000000000000000000b00590000000000000000000000000000000000000000000b00ef1a00000000000000000000000000000000000000000b00fe0500000000000000000000000000000000000000000b00db2500000000000000000000000000000000000000000b00461300000000000000000000000000000000000000000b002c2200000000000000000000000000000000000000000b002d0800000000000000000000000000000000000000000b00934500000000000000000000000000000000000000000b00ca2000000000000000000000000000000000000000000b00cc4600000000000000000000000000000000000000000b00db2000000000000000000000000000000000000000000b00080000000000000000000000000000000000000000000b00760a00000000000000000000000000000000000000000b00e51900000000000000000000000000000000000000000b00270e00000000000000000000000000000000000000000b00524300000000000000000000000000000000000000000b00be1e00000000000000000000000000000000000000000b00790800000000000000000000000000000000000000000b00441900000000000000000000000000000000000000000b00d03d00000000000000000000000000000000000000000b00fd1200000000000000000000000000000000000000000b00242a00000000000000000000000000000000000000000b00d20100000000000000000000000000000000000000000b00a04800000000000000000000000000000000000000000b00394a00000000000000000000000000000000000000000b001f0100000000000000000000000000000000000000000b00331a00000000000000000000000000000000000000000b00cf2f00000000000000000000000000000000000000000b00702600000000000000000000000000000000000000000b00b00b00000000000000000000000000000000000000000b000b4200000000000000000000000000000000000000000b00e22b00000000000000000000000000000000000000000b00dd2f00000000000000000000000000000000000000000b00b60a00000000000000000000000000000000000000000b006b3d00000000000000000000000000000000000000000b00a53c00000000000000000000000000000000000000000b00b92900000000000000000000000000000000000000000b00d63600000000000000000000000000000000000000000b00dc0e00000000000000000000000000000000000000000b00f82900000000000000000000000000000000000000000b00702100000000000000000000000000000000000000000b00b22100000000000000000000000000000000000000000b00513600000000000000000000000000000000000000000b00f73300000000000000000000000000000000000000000b00b02700000000000000000000000000000000000000000b00d54600000000000000000000000000000000000000000b00f60c00000000000000000000000000000000000000000b00082a00000000000000000000000000000000000000000b00fd3300000000000000000000000000000000000000000b00393400000000000000000000000000000000000000000b000a0400000000000000000000000000000000000000000b00473d00000000000000000000000000000000000000000b00bb3000000000000000000000000000000000000000000b00240100000000000000000000000000000000000000000b00460500000000000000000000000000000000000000000b005f4700000000000000000000000000000000000000000b002d4b00000000000000000000000000000000000000000b00674700000000000000000000000000000000000000000b00be2600000000000000000000000000000000000000000b00642c00000000000000000000000000000000000000000b003a3200000000000000000000000000000000000000000b00684500000000000000000000000000000000000000000b00673a00000000000000000000000000000000000000000b00101a00000000000000000000000000000000000000000b00b73100000000000000000000000000000000000000000b005b0e00000000000000000000000000000000000000000b007c2b00000000000000000000000000000000000000000b00441400000000000000000000000000000000000000000b006e4400000000000000000000000000000000000000000b00034700000000000000000000000000000000000000000b00f00c00000000000000000000000000000000000000000b00ec0000000000000000000000000000000000000000000b00df1800000000000000000000000000000000000000000b00f43300000000000000000000000000000000000000000b00e32200000000000000000000000000000000000000000b00d43800000000000000000000000000000000000000000b002e2900000000000000000000000000000000000000000b00464400000000000000000000000000000000000000000b000a2f00000000000000000000000000000000000000000b007f3700000000000000000000000000000000000000000b00624900000000000000000000000000000000000000000b00192a00000000000000000000000000000000000000000b00cc0800000000000000000000000000000000000000000b00330800000000000000000000000000000000000000000b00b43000000000000000000000000000000000000000000b007d0e00000000000000000000000000000000000000000b00370500000000000000000000000000000000000000000b00b44300000000000000000000000000000000000000000b00903a00000000000000000000000000000000000000000b00ba0300000000000000000000000000000000000000000b00334100000000000000000000000000000000000000000b00910600000000000000000000000000000000000000000b00f50d00000000000000000000000000000000000000000b002c3f00000000000000000000000000000000000000000b006c3900000000000000000000000000000000000000000b00662d00000000000000000000000000000000000000000b00f64600000000000000000000000000000000000000000b00664600000000000000000000000000000000000000000b008c4b00000000000000000000000000000000000000000b00e62800000000000000000000000000000000000000000b00cc1500000000000000000000000000000000000000000b00fd2d00000000000000000000000000000000000000000b00113d00000000000000000000000000000000000000000b00e31100000000000000000000000000000000000000000b00450f00000000000000000000000000000000000000000b005f3100000000000000000000000000000000000000000b00243000000000000000000000000000000000000000000b00154200000000000000000000000000000000000000000b00a41900000000000000000000000000000000000000000b00152600000000000000000000000000000000000000000b00fc4400000000000000000000000000000000000000000b00303200000000000000000000000000000000000000000b00c20200000000000000000000000000000000000000000b00d41300000000000000000000000000000000000000000b00ec0400000000000000000000000000000000000000000b00f71100000000000000000000000000000000000000000b00ae4700000000000000000000000000000000000000000b00453200000000000000000000000000000000000000000b00801800000000000000000000000000000000000000000b00cd0600000000000000000000000000000000000000000b00eb3b00000000000000000000000000000000000000000b001a3000000000000000000000000000000000000000000b00bc3e00000000000000000000000000000000000000000b005b0900000000000000000000000000000000000000000b006a2600000000000000000000000000000000000000000b00c01700000000000000000000000000000000000000000b00632200000000000000000000000000000000000000000b00892b00000000000000000000000000000000000000000b00071000000000000000000000000000000000000000000a00f00c00000000000000000000000000000000000000000a00200d00000000000000000000000000000000000000000a00500d00000000000000000000000000000000000000000b008c0600000000000000000000000000000000000000000b00173500000000000000000000000000000000000000000b00db2c00000000000000000000000000000000000000000b00091800000000000000000000000000000000000000000b00121800000000000000000000000000000000000000000b000e2d00000000000000000000000000000000000000000b004c1500000000000000000000000000000000000000000b00b94400000000000000000000000000000000000000000300a84201000000000000000000000000000000000000000300b642010000000000000000000000000000000000000003007877010000000000000000000000000000000000000003007a7701000000000000000000000000000000000000000300bc7801000000000000000000000000000000000000000300a07a01000000000000000000000000000000000000000300f67a010000000000000000000000000000000000000003006e7e010000000000000000000000000000000000000003007c7e01000000000000000000000000000000000000000300fa7f010000000000000000000000000000000000000003000c80010000000000000000000000000000000000000003001e80010000000000000000000000000000000000000003002c80010000000000000000000000000000000000000003003a8001000000000000000000000000000000000000000300488001000000000000000000000000000000000000000300b880010000000000000000000000000000000000000003007482010000000000000000000000000000000000000003002883010000000000000000000000000000000000000003006083010000000000000000000000000000000000000003006a83010000000000000000000000000000000000000003002084010000000000000000000000000000000000000003005a84010000000000000000000000000000000000000003007a8501000000000000000000000000000000000000000300128601000000000000000000000000000000000000000300208601000000000000000000000000000000000000000300368601000000000000000000000000000000000000000300d8860100000000000000000000000000000000000000030048870100000000000000000000000000973800000400f1ff000000000000000000000000000000009d38000000000300eea40100000000000000000000000000a038000000000300bca50100000000000000000000000000a338000000000300e4a90100000000000000000000000000a6380000000003000aaa0100000000000000000000000000a938000000000300baa50100000000000000000000000000ad38000000000300aaa50100000000000000000000000000b138000000000300e0a90100000000000000000000000000b63800000000030098a60100000000000000000000000000bb38000000000300e0a50100000000000000000000000000c03800000000030082a80100000000000000000000000000c538000000000300dca50100000000000000000000000000ca38000000000300aca60100000000000000000000000000cf3800000000030058a60100000000000000000000000000d43800000000030016a60100000000000000000000000000d9380000000003001aa90100000000000000000000000000de3800000000030026a60100000000000000000000000000e3380000000003007ea60100000000000000000000000000e8380000000003008aa60100000000000000000000000000ed380000000003006ca80100000000000000000000000000f23800000000030060a70100000000000000000000000000f7380000000003004aa90100000000000000000000000000fc380000000003008ca801000000000000000000000000000139000000000300f6a601000000000000000000000000000639000000000300faa701000000000000000000000000000b3900000000030042a80100000000000000000000000000103900000000030068a8010000000000000000000000000015390000000003008ea601000000000000000000000000001a39000000000300aea801000000000000000000000000001f3900000000030024a90100000000000000000000000000243900000000030074a901000000000000000000000000002939000000000300f4a501000000000000000000000000002e39000000000300faa901000000000000000000000000003439000000000300fea901000000000000000000000000003a39000000000300e6a901000000000000000000000000004039000000000300eaaa01000000000000000000000000004639000000000300caab01000000000000000000000000004c39000000000300eeaa0100000000000000000000000000523900000000030056ab01000000000000000000000000005839000000000300d0ab01000000000000000000000000005e39000000000300ccab010000000000000000000000000064390000000003006caa01000000000000000000000000006a3900000000030040ab01000000000000000000000000007039000000000300e6ab010000000000000000000000000076390000000003000cab01000000000000000000000000007c3900000000030006ab01000000000000000000000000008239000000000300d6ab010000000000000000000000000088390000000003002aab01000000000000000000000000008e39000000000300eaab010000000000000000000000000094390000000003006eab01000000000000000000000000009a3900000000030068ab0100000000000000000000000000a039000000000300daab0100000000000000000000000000a63900000000030096ab0100000000000000000000000000ac39000000000300b8ab0100000000000000000000000000b239000000000300b6ab0100000000000000000000000000b839000000000300b2ab0100000000000000000000000000be3900000000030020ab0100000000000000000000000000c43900000000030080ab0100000000000000000000000000e039000002020300eea4010000000000ce00000000000000e739000002020300bca50100000000002804000000000000ee39000002020300e4a90100000000002600000000000000f5390000020203000aaa010000000000e601000000000000ca39000012000300ea26010000000000181b000000000000d939000010000300d4260100000000000000000000000000002e726f64617461002e65685f6672616d65002e74657874002e7364617461002e64617461002e627373002e64656275675f616262726576002e64656275675f696e666f002e64656275675f6172616e676573002e64656275675f72616e676573002e64656275675f737472002e64656275675f7075626e616d6573002e64656275675f7075627479706573002e72697363762e61747472696275746573002e64656275675f6c696e65002e636f6d6d656e74002e73796d746162002e7368737472746162002e73747274616200007374616b652e643261633065616565393339383164632d6367752e30002e4c706372656c5f686930005f5a4e37636b625f73746433656e7634415247563137683036373561626564353032343439613545005f5a4e35616c6c6f63377261775f7665633139526177566563244c54245424432441244754243131616c6c6f636174655f696e3137683961373435623837316432623838663945002e4c706372656c5f686931002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e343330002e4c706372656c5f686933002e4c706372656c5f686932005f5a4e34636f726533707472353564726f705f696e5f706c616365244c54246d6f6c6563756c652e2e6572726f722e2e566572696669636174696f6e4572726f72244754243137683936383830623737653965663033383845005f5f727573745f6465616c6c6f63005f5a4e39305f244c54247574696c2e2e6572726f722e2e4572726f72247532302461732475323024636f72652e2e636f6e766572742e2e46726f6d244c5424636b625f7374642e2e6572726f722e2e5379734572726f7224475424244754243466726f6d3137686233643163343538633564356263343545002e4c706372656c5f686934002e4c706372656c5f686935002e4c706372656c5f686936005f5a4e34636f726535736c69636535696e64657837345f244c5424696d706c2475323024636f72652e2e6f70732e2e696e6465782e2e496e646578244c542449244754242475323024666f72247532302424753562245424753564242447542435696e6465783137683064326565363561653136626361336545005f5a4e3131315f244c5424616c6c6f632e2e7665632e2e566563244c54245424475424247532302461732475323024616c6c6f632e2e7665632e2e737065635f66726f6d5f697465725f6e65737465642e2e5370656346726f6d497465724e6573746564244c5424542443244924475424244754243966726f6d5f697465723137683032353562336632346332623633633445005f5a4e35616c6c6f63337665633136566563244c542454244324412447542434707573683137683832346530366138613965323339383745005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f7233616e793137683031323866356465313834336464653445002e4c706372656c5f686938002e4c706372656c5f686937005f5a4e3130325f244c5424636b625f7374616e64616c6f6e655f74797065732e2e67656e6572617465642e2e626c6f636b636861696e2e2e42797465735265616465722475323024617324753230246d6f6c6563756c652e2e7072656c7564652e2e52656164657224475424367665726966793137683135663233383466353032373265326345005f5a4e386d6f6c6563756c6535627974657335427974657335736c6963653137683339643866386561613338343133646245002e4c706372656c5f686939002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e3936002e4c706372656c5f68693130002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e3234005f5a4e386d6f6c6563756c6535627974657335427974657335736c6963653137683133633337653065643765643238336345005f5a4e39385f244c54246d6f6c6563756c65322e2e7265616465722e2e437572736f72247532302461732475323024636f72652e2e636f6e766572742e2e46726f6d244c5424616c6c6f632e2e7665632e2e566563244c542475382447542424475424244754243466726f6d3137686365383937663564613837343036643045005f5a4e396d6f6c6563756c65323672656164657236437572736f723135736c6963655f62795f6f66667365743137683635646335653064333235363034343945005f5a4e396d6f6c6563756c6532367265616465723130385f244c5424696d706c2475323024636f72652e2e636f6e766572742e2e46726f6d244c54246d6f6c6563756c65322e2e7265616465722e2e437572736f72244754242475323024666f722475323024616c6c6f632e2e7665632e2e566563244c5424753824475424244754243466726f6d3137683965653331373661666261663535343545005f5a4e36345f244c5424616c6c6f632e2e72632e2e5263244c54245424475424247532302461732475323024636f72652e2e6f70732e2e64726f702e2e44726f70244754243464726f703137683663346239333364656266363135663545002e4c706372656c5f68693136002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e383436002e4c706372656c5f68693138002e4c706372656c5f68693137002e4c706372656c5f68693139002e4c706372656c5f68693230002e4c706372656c5f68693231002e4c706372656c5f68693233002e4c706372656c5f68693232005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243135636f70795f66726f6d5f736c69636531376c656e5f6d69736d617463685f6661696c3137686531663934356265353831313135613845002e4c706372656c5f68693131007374722e342e3436005f5a4e34636f72653970616e69636b696e673570616e69633137686437373538656430613265383739363145005f5a4e39385f244c5424636b625f7374642e2e686967685f6c6576656c2e2e517565727949746572244c54244624475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137686231366136333531633137303061613745005f5a4e37636b625f7374643130686967685f6c6576656c31346c6f61645f63656c6c5f646174613137686438663961623933373437336639633645005f5a4e396d6f6c6563756c65323672656164657236437572736f7232307461626c655f736c6963655f62795f696e6465783137686232343839353738643638326165663045005f5a4e347574696c3668656c70657231356765745f7363726970745f686173683137683861333134336361336163636135633445005f5a4e37636b625f7374643130686967685f6c6576656c31396c6f61645f63656c6c5f6c6f636b5f686173683137686238376330343133623735373432633545005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f72656164657237547970654964733134787564745f747970655f686173683137686334653636633566343738343237356145005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f726561646572375479706549647331397374616b655f736d745f636f64655f686173683137683939313230643232643561376161363745005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f726561646572375479706549647331377374616b655f736d745f747970655f69643137683133613730383736373561386135323245005f5a4e347574696c3668656c70657232376765745f63656c6c5f636f756e745f62795f747970655f686173683137683636366663636666636434353161366445005f5a4e347574696c3668656c7065723230636865636b5f787564745f747970655f686173683137683036636334386162663931333435343345005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231355374616b65417443656c6c4461746131366d657461646174615f747970655f69643137683136353731366261626264366365656645005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f72656164657237547970654964733138636865636b706f696e745f747970655f69643137683062376537323033303666383865346345005f5a4e347574696c3668656c70657232316765745f787564745f62795f747970655f686173683137686133323939383965653034636166616145002e4c706372656c5f68693238007374722e302e333235002e4c706372656c5f68693132002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3436002e4c706372656c5f68693133002e4c616e6f6e2e65383134633736363361666663333138633766356639363865643531663662352e3139002e4c706372656c5f68693134002e4c706372656c5f68693135005f5a4e34636f726536726573756c743133756e777261705f6661696c65643137683030653934303161326339653536633045005f5a4e347574696c3668656c70657233306765745f7374616b655f61745f646174615f62795f6c6f636b5f686173683137683536356232313136353933333665623945005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231345374616b65496e666f44656c7461313169735f696e6372656173653137683166386136356661303836623163316645005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231355374616b65417443656c6c446174613564656c74613137683762333332613765343438316530613845005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231345374616b65496e666f44656c746136616d6f756e743137683736303137613463316430633135626445005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231345374616b65496e666f44656c74613138696e61756775726174696f6e5f65706f63683137683538323561303933383837366165313345005f5a4e347574696c3668656c70657231376765745f63757272656e745f65706f63683137683433313039626562306665666534313945002e4c706372656c5f68693236002e4c706372656c5f68693237002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3438002e4c706372656c5f68693234002e4c706372656c5f68693235002e4c616e6f6e2e36633237623166666234666234346562313164656530663863336331326232322e32002e4c706372656c5f68693239002e4c706372656c5f68693330002e4c706372656c5f68693331002e4c706372656c5f68693332002e4c706372656c5f68693333002e4c706372656c5f68693334002e4c706372656c5f68693335002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e34002e4c706372656c5f68693336007374722e30002e4c706372656c5f68693337007374722e31002e4c706372656c5f68693430002e4c706372656c5f68693339002e4c706372656c5f6869333800727573745f626567696e5f756e77696e64005f5a4e37636b625f7374643873797363616c6c73366e617469766534657869743137683163616638653234666532613530323145005f5f72675f616c6c6f63005f5a4e3130365f244c542462756464795f616c6c6f632e2e6e6f6e5f746872656164736166655f616c6c6f632e2e4e6f6e54687265616473616665416c6c6f63247532302461732475323024636f72652e2e616c6c6f632e2e676c6f62616c2e2e476c6f62616c416c6c6f632447542435616c6c6f633137683966656332343337626566343266383945005f5f72675f6465616c6c6f63005f5a4e3130365f244c542462756464795f616c6c6f632e2e6e6f6e5f746872656164736166655f616c6c6f632e2e4e6f6e54687265616473616665416c6c6f63247532302461732475323024636f72652e2e616c6c6f632e2e676c6f62616c2e2e476c6f62616c416c6c6f6324475424376465616c6c6f633137686530336235656339643238613732396445005f5f72675f7265616c6c6f63005f5f72675f616c6c6f635f7a65726f6564005f5a4e35616c6c6f63377261775f766563313763617061636974795f6f766572666c6f773137683736396433373734353939336431626545005f5a4e34636f72653970616e69636b696e67313870616e69635f6e6f756e77696e645f666d743137683133386130386530383963323036303445005f5f72646c5f6f6f6d002e4c706372656c5f68693431002e4c706372656c5f68693432002e4c706372656c5f68693433002e4c706372656c5f68693434002e4c706372656c5f68693435002e4c706372656c5f68693436002e4c706372656c5f68693437002e4c706372656c5f68693438005f5a4e396d6f6c6563756c65323672656164657238355f244c5424696d706c2475323024636f72652e2e636f6e766572742e2e46726f6d244c54246d6f6c6563756c65322e2e7265616465722e2e437572736f72244754242475323024666f7224753230247538244754243466726f6d3137686461653235633931336631613435396545002e4c706372656c5f68693439002e4c706372656c5f68693530002e4c706372656c5f68693531002e4c706372656c5f68693532005f5a4e396d6f6c6563756c65323672656164657238365f244c5424696d706c2475323024636f72652e2e636f6e766572742e2e46726f6d244c54246d6f6c6563756c65322e2e7265616465722e2e437572736f72244754242475323024666f722475323024753634244754243466726f6d3137686232663035653938653831303635333145002e4c706372656c5f68693533002e4c706372656c5f68693534002e4c706372656c5f68693535002e4c706372656c5f68693536002e4c706372656c5f68693537002e4c706372656c5f68693538005f5a4e3131626c616b6532625f7265663131626c616b6532625f7265663138626c616b6532625f696e69745f706172616d3137683431613831343963666239633164343445002e4c706372656c5f68693539005f5a4e3131626c616b6532625f7265663131626c616b6532625f7265663130626c616b6532625f49563137686532356438333932346363316638393145005f5a4e3131626c616b6532625f7265663131626c616b6532625f7265663134626c616b6532625f7570646174653137683337646637643338333264666265336545005f5a4e3131626c616b6532625f7265663131626c616b6532625f7265663136626c616b6532625f636f6d70726573733137683531363361326435303733336262323945002e4c43504931395f30002e4c43504931395f31002e4c43504931395f32002e4c43504931395f33002e4c43504931395f34002e4c43504931395f35002e4c43504931395f36002e4c43504931395f37002e4c706372656c5f68693630002e4c706372656c5f68693631002e4c706372656c5f68693632002e4c706372656c5f68693633002e4c706372656c5f68693634002e4c706372656c5f68693635002e4c706372656c5f68693636002e4c706372656c5f68693637005f5a4e313162756464795f616c6c6f63313162756464795f616c6c6f6331304275646479416c6c6f63336e65773137683039343964346234353436656265666245005f5a4e313162756464795f616c6c6f63313162756464795f616c6c6f6337726f756e6475703137686533656266373734346663663366363345002e4c706372656c5f68693735007374722e342e3336005f5a4e313162756464795f616c6c6f63313162756464795f616c6c6f63366e626c6f636b3137683537623963376462363561386133343745005f5a4e313162756464795f616c6c6f63313162756464795f616c6c6f6331304275646479416c6c6f633131626c6f636b5f696e6465783137683333633165376336333564613363643945005f5a4e34636f7265366f7074696f6e31336578706563745f6661696c65643137686332333330616533386638616564396545002e4c706372656c5f68693830002e4c706372656c5f68693736002e4c706372656c5f68693737002e4c706372656c5f68693638002e4c706372656c5f68693730007374722e322e3337002e4c706372656c5f68693731007374722e332e3338002e4c706372656c5f68693732002e4c706372656c5f68693733007374722e312e3335002e4c706372656c5f68693734002e4c706372656c5f68693831002e4c706372656c5f68693738007374722e302e3334002e4c706372656c5f68693639002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3135002e4c706372656c5f68693832002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3238005f5a4e34636f72653970616e69636b696e67313370616e69635f646973706c61793137683538303536323433613031393534316645002e4c706372656c5f68693739002e4c706372656c5f68693833002e4c706372656c5f68693834002e4c706372656c5f68693835002e4c706372656c5f68693836002e4c706372656c5f68693837002e4c706372656c5f68693839002e4c706372656c5f68693930002e4c706372656c5f68693838002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3338005f5a4e313162756464795f616c6c6f633130666173745f616c6c6f633946617374416c6c6f63336e65773137683239303962396561363461333531383845002e4c706372656c5f68693932002e4c706372656c5f68693931002e4c706372656c5f68693933002e4c706372656c5f68693934005f5a4e357374616b6535414c4c4f433137683735313734646435353830643734633445002e4c706372656c5f68693938002e4c706372656c5f6869313033002e4c706372656c5f6869313034002e4c706372656c5f6869313031002e4c706372656c5f6869313035002e4c706372656c5f6869313036002e4c706372656c5f6869313032002e4c706372656c5f68693937002e4c706372656c5f68693939002e4c706372656c5f6869313030002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e32002e4c706372656c5f68693935002e4c706372656c5f68693936002e4c706372656c5f6869313037002e4c706372656c5f6869313038002e4c706372656c5f6869313039002e4c706372656c5f6869313133002e4c706372656c5f6869313132002e4c706372656c5f6869313136002e4c706372656c5f6869313138002e4c706372656c5f6869313139002e4c706372656c5f6869313230002e4c706372656c5f6869313137002e4c706372656c5f6869313130002e4c706372656c5f6869313131002e4c706372656c5f6869313134002e4c706372656c5f6869313135005f5a4e35616c6c6f63377261775f7665633139526177566563244c54245424432441244754243131616c6c6f636174655f696e3137683334393639363464643031633234363645005f5a4e35616c6c6f63377261775f7665633139526177566563244c542454244324412447542437726573657276653231646f5f726573657276655f616e645f68616e646c653137686234636364626536643135363830353445002e4c706372656c5f6869313231007374722e302e3434005f5f727573745f616c6c6f63005f5f727573745f616c6c6f635f6572726f725f68616e646c6572005f5a4e35616c6c6f63377261775f7665633139526177566563244c5424542443244124475424313467726f775f616d6f7274697a65643137683131313435313531653037646531613245005f5a4e35616c6c6f63377261775f766563313166696e6973685f67726f773137683362363537323731663362336132663345005f5a4e35616c6c6f63377261775f7665633139526177566563244c54245424432441244754243136726573657276655f666f725f707573683137683364383734353931323332303230376445002e4c706372656c5f6869313232002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e313734002e4c706372656c5f6869313233002e4c706372656c5f6869313234005f5a4e36315f244c5424636b625f7374642e2e6572726f722e2e5379734572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683863383033303266623836336136303845002e4c706372656c5f6869313235002e4c4a544933395f30002e4c424233395f31002e4c706372656c5f6869313236002e4c616e6f6e2e34313466363731613135666237623063306532636261396133343630323939342e3339002e4c424233395f32002e4c706372656c5f6869313237002e4c616e6f6e2e34313466363731613135666237623063306532636261396133343630323939342e3338002e4c424233395f33002e4c706372656c5f6869313238002e4c616e6f6e2e34313466363731613135666237623063306532636261396133343630323939342e3336002e4c706372656c5f6869313239002e4c616e6f6e2e34313466363731613135666237623063306532636261396133343630323939342e3337002e4c424233395f34002e4c706372656c5f6869313330002e4c424233395f36002e4c706372656c5f6869313331002e4c616e6f6e2e34313466363731613135666237623063306532636261396133343630323939342e3333002e4c706372656c5f6869313332002e4c616e6f6e2e34313466363731613135666237623063306532636261396133343630323939342e3334005f5a4e34636f726533666d7439466f726d6174746572323564656275675f7475706c655f6669656c64315f66696e6973683137683963326264643732306464613133376545005f5a4e34636f726533707472323864726f705f696e5f706c616365244c542424524624753634244754243137683536663832373834643464373061633345005f5a4e37636b625f7374643130686967685f6c6576656c31396c6f61645f63656c6c5f747970655f686173683137686661353738353337303831333261613945005f5a4e34636f7265336f70733866756e6374696f6e36466e4f6e63653963616c6c5f6f6e63653137683331326365396462383432326365623645005f5a4e34636f72653370747231303264726f705f696e5f706c616365244c542424524624636f72652e2e697465722e2e61646170746572732e2e636f706965642e2e436f70696564244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c542475382447542424475424244754243137683465633534623435323134663763393045002e4c43504934385f30005f5a4e34636f726533666d74336e756d33696d7037666d745f7536343137683238366534643532373433386334363745002e4c706372656c5f6869313333002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333234002e4c706372656c5f6869313334002e4c706372656c5f6869313335002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3233005f5a4e34636f726533666d7439466f726d617474657231327061645f696e74656772616c3137686238656639343965396131613633346545005f5a4e34636f726533666d7439466f726d617474657231327061645f696e74656772616c313277726974655f7072656669783137683834663538656430383761336264393345002e4c43504935315f30002e4c43504935315f31005f5a4e34636f726533666d7439466f726d6174746572337061643137683433336537613934646232626438653245002e4c706372656c5f6869313336002e4c706372656c5f6869313337005f5a4e34636f726533666d743577726974653137683537653362636463656237646630393145002e4c706372656c5f6869313338005f5a4e36305f244c5424636f72652e2e63656c6c2e2e426f72726f774572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137686163386261333334363731373261333845002e4c706372656c5f6869313339002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e313730005f5a4e36335f244c5424636f72652e2e63656c6c2e2e426f72726f774d75744572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683636336332373865383138373636393045002e4c706372656c5f6869313430002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e313731005f5a4e34636f726533666d74336e756d35335f244c5424696d706c2475323024636f72652e2e666d742e2e4c6f7765724865782475323024666f7224753230246936342447542433666d743137686632356530653835343735353364373145002e4c706372656c5f6869313431002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333232002e4c43504936305f30002e4c43504936305f31002e4c43504936305f32005f5a4e36385f244c5424636f72652e2e666d742e2e6275696c646572732e2e50616441646170746572247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f7374723137686539366438303337316562386433343445002e4c706372656c5f6869313432002e4c706372656c5f6869313433002e4c706372656c5f6869313434002e4c706372656c5f6869313435005f5a4e34636f726533666d74355772697465313077726974655f636861723137686664666234386663643336373461323845005f5a4e34636f726533666d743557726974653977726974655f666d743137683364623431343565346436363932376245002e4c706372656c5f6869313436002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333237005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f7374723137683865303931326361326264646233386345005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e577269746524475424313077726974655f636861723137683239666437616639333939643762333645005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f666d743137683565373464633863623261616161323645002e4c706372656c5f6869313437005f5a4e34636f726533666d74386275696c64657273313044656275675475706c65356669656c643137686134393061356537663734366534656245002e4c706372656c5f6869313439002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e323933002e4c706372656c5f6869313530002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333030002e4c706372656c5f6869313438002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333031002e4c706372656c5f6869313531002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e323839002e4c706372656c5f6869313532002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e323932002e4c706372656c5f6869313534002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333032002e4c706372656c5f6869313533002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e313537005f5a4e34325f244c54242452462454247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137686332303631326561373836393861653445002e4c706372656c5f6869313535002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333337005f5a4e36375f244c5424636f72652e2e61727261792e2e54727946726f6d536c6963654572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683532646436363362353834636335356645002e4c706372656c5f6869313536002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e353537002e4c706372656c5f6869313537002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e353333002e4c706372656c5f6869313539002e4c706372656c5f6869313538005f5a4e34636f726533666d74336e756d35335f244c5424696d706c2475323024636f72652e2e666d742e2e55707065724865782475323024666f7224753230246936342447542433666d743137683464336136353331313038303933376445002e4c706372656c5f6869313630005f5a4e3133325f244c5424616c6c6f632e2e7665632e2e566563244c5424542443244124475424247532302461732475323024616c6c6f632e2e7665632e2e737065635f657874656e642e2e53706563457874656e64244c54242452462454244324636f72652e2e736c6963652e2e697465722e2e49746572244c5424542447542424475424244754243131737065635f657874656e643137683464663561353366366631653763336445005f5a4e35616c6c6f63377261775f7665633139526177566563244c542454244324412447542437726573657276653231646f5f726573657276655f616e645f68616e646c653137686332663335393562613638613033633645005f5f727573745f7265616c6c6f63005f5a4e34325f244c54242452462454247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683431323134373832613466363464656645005f5f727573745f616c6c6f635f7a65726f6564005f5a4e35616c6c6f63337665633136566563244c54245424432441244754243131657874656e645f776974683137683935323361376565386561616133316645005f5a4e35616c6c6f63377261775f7665633139526177566563244c542454244324412447542437726573657276653231646f5f726573657276655f616e645f68616e646c653137686534386235666233366361343936633545005f5a4e35616c6c6f63377261775f766563313166696e6973685f67726f773137686465323762646133633136313431313345005f5a4e396d6f6c6563756c65323672656164657237726561645f61743137686436323832346538376630396538383045002e4c706372656c5f6869313730007374722e312e323830002e4c706372656c5f6869313633002e4c706372656c5f6869313634002e4c706372656c5f6869313631002e4c706372656c5f6869313632002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e31002e4c706372656c5f6869313639002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3136002e4c706372656c5f6869313731002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3139002e4c706372656c5f6869313635002e4c706372656c5f6869313636002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e36002e4c706372656c5f6869313637002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3132002e4c706372656c5f6869313638002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3134005f5a4e36315f244c54246d6f6c6563756c65322e2e7265616465722e2e4572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683238346238363235356264316239336545002e4c706372656c5f6869313732002e4c7377697463682e7461626c652e5f5a4e36315f244c54246d6f6c6563756c65322e2e7265616465722e2e4572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683238346238363235356264316239336545002e4c706372656c5f6869313733002e4c7377697463682e7461626c652e5f5a4e36315f244c54246d6f6c6563756c65322e2e7265616465722e2e4572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d7431376832383462383632353562643162393365452e333731005f5a4e396d6f6c6563756c65323672656164657236437572736f723876616c69646174653137683930306131623931383065653939313845002e4c706372656c5f6869313736002e4c706372656c5f6869313734002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e32002e4c706372656c5f6869313735002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e33002e4c706372656c5f6869313737002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3238005f5a4e396d6f6c6563756c65323672656164657236437572736f723133756e7061636b5f6e756d6265723137683635326430373132666263326536343145002e4c706372656c5f6869313738002e4c706372656c5f6869313739002e4c706372656c5f6869313830002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3331002e4c706372656c5f6869313831002e4c706372656c5f6869313839002e4c706372656c5f6869313832002e4c706372656c5f6869313833002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3335002e4c706372656c5f6869313834002e4c706372656c5f6869313838002e4c706372656c5f6869313835002e4c706372656c5f6869313836002e4c706372656c5f6869313837002e4c706372656c5f6869313930002e4c706372656c5f6869313931002e4c706372656c5f6869313932002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3430002e4c706372656c5f6869313933002e4c706372656c5f6869313934002e4c706372656c5f6869313935002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3538002e4c706372656c5f6869313936002e4c706372656c5f6869313937002e4c706372656c5f6869313938002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3634005f5a4e36395f244c5424616c6c6f632e2e7665632e2e566563244c54247538244754242475323024617324753230246d6f6c6563756c65322e2e7265616465722e2e526561642447542434726561643137683538323363346134366134643066373445002e4c706372656c5f6869313939002e4c706372656c5f6869323030002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3638005f5a4e34636f726533707472343664726f705f696e5f706c616365244c5424616c6c6f632e2e7665632e2e566563244c5424753824475424244754243137683139303635656264313265376238616645002e4c706372656c5f6869323031005f5a4e3130325f244c5424636f72652e2e697465722e2e61646170746572732e2e6d61702e2e4d6170244c5424492443244624475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424387472795f666f6c643137686134643535656336343238393364643045002e4c706372656c5f6869323035002e4c706372656c5f6869323034002e4c706372656c5f6869323032002e4c706372656c5f6869323033002e4c706372656c5f6869323036002e4c4a54493130305f30002e4c42423130305f31002e4c42423130305f32002e4c42423130305f33002e4c42423130305f34002e4c42423130305f35002e4c706372656c5f6869323134002e4c706372656c5f6869323039007374722e322e3433002e4c706372656c5f6869323130002e4c706372656c5f6869323131002e4c706372656c5f6869323132002e4c706372656c5f6869323133002e4c706372656c5f6869323037002e4c706372656c5f6869323038002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3437002e4c706372656c5f6869323136002e4c706372656c5f6869323135002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e313134002e4c706372656c5f6869323137002e4c706372656c5f6869323138002e4c706372656c5f6869323139002e4c706372656c5f6869323230002e4c706372656c5f6869323231002e4c706372656c5f6869323232002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e313139002e4c706372656c5f6869323233005f5a4e357374616b6531315f42554444595f484541503137683862313032653565633363313635316445005f5a4e357374616b6531375f46495845445f424c4f434b5f484541503137686132366633373037356664663339316245002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3134002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3237002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3732002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3733002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3734002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3735002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3736002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3737002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3738002e4c6c696e655f7461626c655f737461727430002e4c6c696e655f7461626c655f737461727431006c69622e63002478002478002478002478002e4c32002e4c33002e4c3335002e4c3437002e4c3132002e4c3739002e4c3830002e4c3134002e4c3135002e4c3136002e4c3831002e4c3138002e4c3230002e4c3231002e4c3738002e4c3235002e4c3236002e4c3237002e4c3238002e4c3331002e4c3332002e4c3333002e4c3334002e4c3330002e4c3137002e4c3239002e4c3130002e4c313433002e4c313437002e4c313438002e4c313439002e4c323033002e4c313532002e4c323034002e4c313735002e4c313736002e4c313632002e4c323031002e4c313737002e4c313638002e4c313730002e4c313738002e4c313731002e4c313733002e4c313536002e4c313539002e4c313630002e4c313631002e4c313634002e4c323035002e4c313537002e4c313637002e4c313534005f5f636b625f7374645f6d61696e005f7374617274006d656d736574006d656d637079006d656d636d70006d656d6d6f7665000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000120000000000000060010100000000006001000000000000680900000000000000000000000000001000000000000000000000000000000009000000010000000200000000000000c80a010000000000c80a0000000000000c0c00000000000000000000000000000800000000000000000000000000000013000000010000000600000000000000d426010000000000d4160000000000001c8500000000000000000000000000000400000000000000000000000000000019000000010000000300000000000000f0bb010000000000f09b00000000000070000000000000000000000000000000080000000000000000000000000000002000000001000000030000000000000060bc010000000000609c000000000000b8000000000000000000000000000000080000000000000000000000000000002600000008000000030000000000000018bd010000000000189d00000000000000200800000000000000000000000000010000000000000000000000000000002b0000000100000000000000000000000000000000000000189d0000000000002802000000000000000000000000000001000000000000000000000000000000390000000100000000000000000000000000000000000000409f0000000000003f230000000000000000000000000000010000000000000000000000000000004500000001000000000000000000000000000000000000007fc200000000000000020000000000000000000000000000010000000000000000000000000000005400000001000000000000000000000000000000000000007fc40000000000005010000000000000000000000000000001000000000000000000000000000000620000000100000030000000000000000000000000000000cfd40000000000005a4c0000000000000000000000000000010000000000000001000000000000006d00000001000000000000000000000000000000000000002921010000000000481b0000000000000000000000000000010000000000000000000000000000007d0000000100000000000000000000000000000000000000713c01000000000024000000000000000000000000000000010000000000000000000000000000008d0000000300007000000000000000000000000000000000953c0100000000002b000000000000000000000000000000010000000000000000000000000000009f0000000100000000000000000000000000000000000000c03c010000000000791c000000000000000000000000000001000000000000000000000000000000ab000000010000003000000000000000000000000000000039590100000000002300000000000000000000000000000001000000000000000100000000000000b400000002000000000000000000000000000000000000006059010000000000f8e2000000000000130000007309000008000000000000001800000000000000bc0000000300000000000000000000000000000000000000583c020000000000ce00000000000000000000000000000001000000000000000000000000000000c60000000300000000000000000000000000000000000000263d020000000000fd39000000000000000000000000000001000000000000000000000000000000",
        "0x7f454c460201010000000000000000000200f3000100000074360100000000004000000000000000c00f04000000000001000000400038000500400016001400060000000400000040000000000000004000010000000000400001000000000018010000000000001801000000000000080000000000000001000000040000000000000000000000000001000000000000000100000000007426000000000000742600000000000000100000000000000100000005000000742600000000000074360100000000007436010000000000be82010000000000be820100000000000010000000000000010000000600000038a901000000000038c902000000000038c902000000000068010000000000006821080000000000001000000000000051e574640600000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000005ca90100000000006ea901000000000080a901000000000098a9010000000000aea9010000000000383802000000000036380200000000003a380200000000003e38020000000000423802000000000056880200000000000093020000000000009302000000000000930200000000002a8a020000000000009302000000000000930200000000008e8c0200000000004a8e0200000000009a8e020000000000617474656d707420746f206164642077697468206f766572666c6f7700000000ee3601000000000018000000000000000800000000000000c8c6010000000000d8a901000000000000000000000000000100000000000000d0c3010000000000d8a9010000000000010000000000000001000000000000005eca010000000000617474656d707420746f206164642077697468206f766572666c6f770000000008c9bcf367e6096a3ba7ca8485ae67bb2bf894fe72f36e3cf1361d5f3af54fa5d182e6ad7f520e511f6c3e2b8c68059b6bbd41fbabd9831f79217e1319cde05bd8a901000000000000000000000000000100000000000000c2bb010000000000617474656d707420746f207368696674206c6566742077697468206f766572666c6f7700000000000000000000000000617474656d707420746f206d756c7469706c792077697468206f766572666c6f77000000000000000000000000000000617474656d707420746f2073756274726163742077697468206f766572666c6f77000000000000000000000000000000617474656d707420746f2073686966742072696768742077697468206f766572666c6f77000000000000000000000000617474656d707420746f206164642077697468206f766572666c6f776c6561662073697a65206d75737420626520616c69676e20746f20313620627974657300dc0301000000000023000000000000007265717569726573206d6f7265206d656d6f727920737061636520746f20696e697469616c697a65204275646479416c6c6f630000000000100401000000000033000000000000006f7574206f66206d656d6f72790000000000000000000000617474656d707420746f20646976696465206279207a65726f00000000000000617474656d707420746f206164642077697468206f766572666c6f77427974655265616465724279746533325265616465724279746573526561646572000000617474656d707420746f2073756274726163742077697468206f766572666c6f7753637269707452656164657243656c6c496e7075745265616465725769746e65737341726773526561646572556e6b6e6f776e00000000d8a9010000000000080000000000000008000000000000004ac6010000000000456e636f64696e674f766572666c6f7776616c69646174654c656e6774684e6f74456e6f75676800d8a9010000000000080000000000000008000000000000004ac60100000000004974656d4d697373696e67496e6465784f75744f66426f756e64000000000000617474656d707420746f206164642077697468206f766572666c6f7729426f72726f774572726f72426f72726f774d75744572726f725b002eb3010000000000180000000000000008000000000000006ebc0100000000002abe010000000000debe0100000000002020202052656164446174612c0a2c20280a282c0a5d307830303031303230333034303530363037303830393130313131323133313431353136313731383139323032313232323332343235323632373238323933303331333233333334333533363337333833393430343134323433343434353436343734383439353035313532353335343535353635373538353936303631363236333634363536363637363836393730373137323733373437353736373737383739383038313832383338343835383638373838383939303931393239333934393539363937393839392eb30100000000000800000000000000080000000000000016bf01000000000020bf010000000000d6bf01000000000028290000000000002eb301000000000008000000000000000800000000000000bac301000000000054727946726f6d536c6963654572726f72636b622d64656661756c742d68617368616c726561647920626f72726f77656400000000000000d8a901000000000000000000000000000100000000000000c2bb010000000000616c7265616479206d757461626c7920626f72726f776564d8a901000000000000000000000000000100000000000000b0bb010000000000d8a9010000000000010000000000000001000000000000005eca010000000000617474656d707420746f206164642077697468206f766572666c6f77726561645f6174206069662073697a65203c20726561645f6c656e60726561645f6174206069662064732e63616368655f73697a65203e2064732e6d61785f63616368655f73697a6560726561645f617420606966206375722e6f6666736574203c2064732e73746172745f706f696e74207c7c202e2e2e60726561645f61742060696620726561645f706f696e74202b20726561645f6c656e203e2064732e63616368655f73697a656076616c69646174653a2073697a65203e206375722e736f757263652e746f74616c5f73697a65756e7061636b5f6e756d6265726765745f6974656d5f636f756e74636f6e766572745f746f5f753634636f6e766572745f746f5f753136636f6e766572745f746f5f7538636f6e7665727420746f205665633c75383e000000000016d001000000000018000000000000000800000000000000e2ce0100000000004669656c64436f756e744f75744f66426f756e64556e6b6e6f776e4974656d4f6666736574486561646572546f74616c53697a65436f6d6d6f6e617373657274696f6e206661696c65643a20696478203c204341504143495459000000000000000000000000000000000000000000000000000000000000000063616c6c656420604f7074696f6e3a3a756e77726170282960206f6e206120604e6f6e65602076616c7565000000617474656d707420746f206164642077697468206f766572666c6f7700000000617373657274696f6e206661696c65643a206f666673657420213d2030202626206f6666736574203c3d206c656e63616c6c65642060526573756c743a3a756e77726170282960206f6e20616e2060457272602076616c756500000000000000d8a901000000000000000000000000000100000000000000d0c3010000000000d8a90100000000001000000000000000080000000000000046a9010000000000ee3601000000000018000000000000000800000000000000c8c6010000000000617373657274696f6e206661696c65643a20656467652e686569676874203d3d2073656c662e686569676874202d2031617373657274696f6e206661696c65643a2073656c662e686569676874203e2030617373657274696f6e206661696c65643a207372632e6c656e2829203d3d206473742e6c656e2829617373657274696f6e206661696c65643a20656467652e686569676874203d3d2073656c662e6e6f64652e686569676874202d2031617373657274696f6e206661696c65643a20636f756e74203e2030617373657274696f6e206661696c65643a206f6c645f72696768745f6c656e202b20636f756e74203c3d204341504143495459617373657274696f6e206661696c65643a206f6c645f6c6566745f6c656e203e3d20636f756e74696e7465726e616c206572726f723a20656e746572656420756e726561636861626c6520636f6465617373657274696f6e206661696c65643a206f6c645f6c6566745f6c656e202b20636f756e74203c3d204341504143495459617373657274696f6e206661696c65643a206f6c645f72696768745f6c656e203e3d20636f756e74617373657274696f6e206661696c65643a206d6174636820747261636b5f656467655f696478207b5c6e202020204c6566744f7252696768743a3a4c6566742869647829203d3e20696478203c3d206f6c645f6c6566745f6c656e2c5c6e202020204c6566744f7252696768743a3a52696768742869647829203d3e20696478203c3d2072696768745f6c656e2c5c6e7d617373657274696f6e206661696c65643a206e65775f6c6566745f6c656e203c3d204341504143495459617373657274696f6e206661696c65643a20636865636b706f696e745f646174612e69735f6e6f6e652829617373657274696f6e206661696c65643a207374616b655f61745f646174612e69735f6e6f6e652829617373657274696f6e206661696c65643a2077697468647261775f61745f646174612e69735f6e6f6e65282906000000000000000900000000000000060000000000000006000000000000000b000000000000000a000000000000000a000000000000000400000000000000080000000000000004000000000000009c0901000000000093090100000000008d0901000000000087090100000000007c0901000000000072090100000000006809010000000000200601000000000050050100000000001c0601000000000008c9bcf367e6096a2bf894fe72f36e3c1f6c3e2b8c68059b3ba7ca8485ae67bb79217e1319cde05bd182e6ad7f520e51f1361d5f3af54fa56bbd41fbabd9831f1000000000000000017a5200017801011b0c02001c00000018000000be2700006400000000420e2048810188028903920400000010000000380000000228000010000000000000001c0000004c000000fe270000ee00000000420e304a81018802890392049305002c0000006c000000cc280000d404000000420e80035a810188028903920493059406950796089709980a990b9a0c9b0d100000009c000000702d000068000000000e000028000000b0000000c42d0000dc00000000420e6056810188028903920493059406950796089709980a990b0014000000dc000000742e00003000000000420e104281010014000000f40000008c2e00003000000000420e10428101002c0000000c010000a42e00007a01000000420e900158810188028903920493059406950796089709980a990b9a0c00002c0000003c010000ee2f0000aa01000000420ea0015a810188028903920493059406950796089709980a990b9a0c9b0d2c0000006c01000068310000c001000000420ed0015a810188028903920493059406950796089709980a990b9a0c9b0d2c0000009c010000f83200008201000000420eb0015a810188028903920493059406950796089709980a990b9a0c9b0d2c000000cc0100004a3400005002000000420ed0035a810188028903920493059406950796089709980a990b9a0c9b0d2c000000fc0100006a360000c600000000420e6058810188028903920493059406950796089709980a990b9a0c000000300000002c020000003700009025000000440ef00f74810188028903920493059406950796089709980a990b9a0c9b0d420e801210000000600200005c5c00000a000000000e00001000000074020000525c000008000000000000001000000088020000465c000008000000000000001c0000009c0200003a5c00004e00000000420e304a810188028903920493050018000000bc020000685c00003000000000420e20468101880289030010000000d80200007c5c0000080000000000000010000000ec020000705c000008000000000000001000000000030000645c000008000000000000001000000014030000585c0000080000000000000010000000280300004c5c00000a000000000e0000140000003c030000425c00000e00000000420e10428101001400000054030000385c00000e00000000420e1042810100180000006c0300002e5c00005800000000420e40448101880200000018000000880300006a5c00005800000000420e40448101880200000018000000a4030000a65c00005800000000420e40448101880200000018000000c0030000e25c00005800000000420e40448101880200000018000000dc0300001e5d00005800000000420e40448101880200000018000000f80300005a5d00005800000000420e4044810188020000001800000014040000965d00005800000000420e4044810188020000001800000030040000d25d00005800000000420e404481018802000000140000004c0400000e5e00005200000000420e40428101001800000064040000485e00005800000000420e4044810188020000001400000080040000845e00005200000000420e40428101001800000098040000be5e00004e00000000420e30448101880200000018000000b4040000f05e00005800000000420e40448101880200000018000000d00400002c5f00005800000000420e40448101880200000018000000ec040000685f00008600000000420e3046810188028903001800000008050000d25f00004c00000000420e3044810188020000001800000024050000026000004e00000000420e3044810188020000001800000040050000346000009400000000420e604481018802000000180000005c050000ac6000009400000000420e6044810188020000001c0000007805000024610000bc00000000420ee00348810188028903920400001c00000098050000c06100009a00000000420e2048810188028903920400000020000000b80500003a620000dc00000000440e304c8101880289039204930594060000002c000000dc050000f2620000ee1a000000420ef0035a810188028903920493059406950796089709980a990b9a0c9b0d1c0000000c060000b07d0000f000000000420e60488101880289039204000000180000002c060000807e00007c00000000420e9003468101880289032c00000048060000e07e00001404000000420e80015a810188028903920493059406950796089709980a990b9a0c9b0d1000000078060000c48200003c000000000e0000100000008c060000ec8200000a000000000e000010000000a0060000e28200004c000000000e000010000000b40600001a8300004c000000000e000010000000c806000052830000f4000000000e00002c000000dc06000032840000d403000000420eb00158810188028903920493059406950796089709980a990b9a0c00002c0000000c070000d6870000f203000000420ec0015a810188028903920493059406950796089709980a990b9a0c9b0d200000003c070000988b0000d600000000420e504e81018802890392049305940695070018000000600700004a8c00005200000000420e204681018802890300140000007c070000808c00003400000000420e104281010018000000940700009c8c00007400000000420e50468101880289030014000000b0070000f48c00003600000000420e104281010020000000c8070000128d00006c00000000420e304c81018802890392049305940600000010000000ec0700005a8d000022000000000e00001800000000080000688d00003a00000000420e204681018802890300200000001c080000868d0000fc00000000420e404e81018802890392049305940695070010000000400800005e8e000042000000000e000020000000540800008c8e00005000000000420e304c8101880289039204930594060000001c00000078080000b88e00007400000000420e4048810188028903920400000020000000980800000c8f00006400000000420e304c8101880289039204930594060000001c000000bc0800004c8f00008200000000420e2048810188028903920400000028000000dc080000ae8f00009601000000420e900154810188028903920493059406950796089709980a000010000000080900001891000072000000000e0000140000001c090000769100009200000000420e10428101001000000034090000f091000002000000000000001000000048090000de9100003600000000000000240000005c09000000920000c001000000440ee008648101880289039204930594069507960897091800000084090000989300007a00000000420e40448101880200000018000000a0090000f69300008200000000420e40448101880200000024000000bc0900005c9400006001000000440ee008648101880289039204930594069507960897092c000000e409000094950000c204000000440e800970810188028903920493059406950796089709980a990b9a0c000010000000140a0000269a000018000000000e000010000000280a00002a9a00002400000000420e10100000003c0a00003a9a0000040000000000000010000000500a00002a9a0000020000000000000014000000640a0000189a00004201000000420e30428101002c0000007c0a0000429b0000e401000000420e705a810188028903920493059406950796089709980a990b9a0c9b0d001c000000ac0a0000f69c00005600000000420e304a810188028903920493050024000000cc0a00002c9d00007803000000420e50528101880289039204930594069507960897090014000000f40a00007ca000000e00000000420e1042810100240000000c0b000072a000007e01000000420e80015081018802890392049305940695079608000010000000340b0000c8a10000120000000000000010000000480b0000c6a100001200000000000000140000005c0b0000c4a100000e00000000420e104281010014000000740b0000baa100000e00000000420e1042810100140000008c0b0000b0a100000e00000000420e104281010014000000a40b0000a6a100007000000000420e90014281012c000000bc0b0000fea10000bc01000000420e90015a810188028903920493059406950796089709980a990b9a0c9b0d14000000ec0b00008aa30000b400000000420e104281010014000000040c000026a400003800000000420e4042810100100000001c0c000046a400000a0000000000000014000000300c00003ca40000b600000000420e104281010014000000480c0000daa400003a00000000420e404281010020000000600c0000fca400002001000000420ea0014e810188028903920493059406950720000000840c0000f8a500000001000000420ea0014e81018802890392049305940695071c000000a80c0000d4a600009800000000420e4048810188028903920400000014000000c80c00004ca700000e00000000420e104281010014000000e00c000042a700007200000000420e900142810114000000f80c00009ca700007200000000420e900142810110000000100d0000f6a70000160000000000000018000000240d0000f8a70000a200000000420e40468101880289030014000000400d00007ea800007000000000420e90014281011c000000580d0000d6a800005200000000420e304a810188028903920493050018000000780d000008a900007e00000000420e5046810188028903001c000000940d00006aa900006200000000420e2048810188028903920400000010000000b40d0000aca90000360000000000000010000000c80d0000cea90000300000000000000018000000dc0d0000eaa900004e00000000420e10448101880200000020000000f80d00001caa00008600000000420e504c8101880289039204930594060000001c0000001c0e00007eaa00006800000000420e304a8101880289039204930500180000003c0e0000c6aa00007e00000000420e50468101880289030018000000580e000028ab00005200000000420e20468101880289030018000000740e00005eab00005600000000420e10448101880200000020000000900e000098ab00008201000000420e504e81018802890392049305940695070010000000b40e0000f6ac0000280000000000000010000000c80e00000aad00006200000000420e1018000000dc0e000058ad00006800000000420e30448101880200000014000000f80e0000a4ad00003000000000420e104281010024000000100f0000bcad00006601000000420e80015281018802890392049305940695079608970918000000380f0000faae00006400000000420e30448101880200000018000000540f000042af00007800000000420e40468101880289030018000000700f00009eaf00007e00000000420e4046810188028903001c0000008c0f000000b00000a200000000420e5048810188028903920400000018000000ac0f000082b000007a00000000420e20468101880289030020000000c80f0000e0b00000ba00000000420e504c81018802890392049305940600000010000000ec0f000076b1000010000000000000001c0000000010000072b100008c00000000420e404881018802890392040000001000000020100000deb100004a000000000000001c0000003410000014b200007200000000420e50488101880289039204000000100000005410000066b20000c0000000000e0000140000006810000012b300002800000000420e1042810100140000008010000022b300002800000000420e10428101002c0000009810000032b300001401000000420e6058810188028903920493059406950796089709980a990b9a0c00000010000000c810000016b400006c000000000000002c000000dc1000006eb400007e03000000420ed0035a810188028903920493059406950796089709980a990b9a0c9b0d2c0000000c110000bcb700000603000000420ec0015a810188028903920493059406950796089709980a990b9a0c9b0d2c0000003c11000092ba0000e802000000420ec0015a810188028903920493059406950796089709980a990b9a0c9b0d2c0000006c1100004abd0000d002000000420eb0015a810188028903920493059406950796089709980a990b9a0c9b0d2c0000009c110000eabf0000ae02000000420ea0015a810188028903920493059406950796089709980a990b9a0c9b0d14000000cc11000068c200002800000000420e104281010014000000e411000078c200002800000000420e104281010028000000fc11000088c200002801000000420e6056810188028903920493059406950796089709980a990b00200000002812000084c300006800000000420e404e8101880289039204930594069507002c0000004c120000c8c300000403000000440ea00674810188028903920493059406950796089709980a990b9a0c9b0d100000007c1200009cc6000066000000000e00002c00000090120000eec60000c602000000440ef00474810188028903920493059406950796089709980a990b9a0c9b0d2c000000c012000084c900004602000000420eb0025a810188028903920493059406950796089709980a990b9a0c9b0d2c000000f01200009acb00008e02000000440ef00474810188028903920493059406950796089709980a990b9a0c9b0d2c00000020130000f8cd00000202000000420e90025a810188028903920493059406950796089709980a990b9a0c9b0d2c00000050130000cacf00003629000000440ec0046a810188028903920493059406950796089709980a990b9a0c9b0d1800000080130000d0f800008e00000000420e504681018802890300200000009c13000042f90000cc01000000440ec0045881018802890392049305940600001c000000c0130000eafa0000f600000000440ec004548101880289039204930520000000e0130000c0fb00005402000000440ee0045881018802890392049305940600002800000004140000f0fd00000604000000420ee00156810188028903920493059406950796089709980a990b2c00000030140000ca010100e809000000420ec00158810188028903920493059406950796089709980a990b9a0c00002400000060140000820b01005001000000420e9001528101880289039204930594069507960897092c00000088140000aa0c01000c03000000420ed0015a810188028903920493059406950796089709980a990b9a0c9b0d24000000b8140000860f0100c803000000420ec001508101880289039204930594069507960800001c000000e0140000261301006a00000000420ea00348810188028903920400001800000000150000701301008e00000000420e5046810188028903001c0000001c150000e21301007200000000420e50488101880289039204000000100000003c1500003414010028000000000e00001000000050150000481401001c00000000000000200000006415000050140100da00000000440ed0055881018802890392049305940600002000000088150000061501002a02000000420ec0014c810188028903920493059406000018000000ac1500000c1701003200000000420e10448101880200000028000000c8150000221701001803000000420eb00256810188028903920493059406950796089709980a990b2c000000f41500000e1a01008c03000000420ef0025a810188028903920493059406950796089709980a990b9a0c9b0d2c000000241600006a1d01009003000000420e80035a810188028903920493059406950796089709980a990b9a0c9b0d2c00000054160000ca2001004e04000000420e80035a810188028903920493059406950796089709980a990b9a0c9b0d2000000084160000e82401008601000000420e90014c81018802890392049305940600002c000000a81600004a2601005602000000420ef0015a810188028903920493059406950796089709980a990b9a0c9b0d1c000000d8160000702801009a00000000420e6048810188028903920400000018000000f8160000ea2801007801000000420ea001468101880289032c00000014170000462a01005402000000420ef0015a810188028903920493059406950796089709980a990b9a0c9b0d2c000000441700006a2c01007207000000440ea00674810188028903920493059406950796089709980a990b9a0c9b0d1800000074170000ac3301007400000000440eb0044c8101880289033000000090170000043401004a3a000000440ef00f74810188028903920493059406950796089709980a990b9a0c9b0d420e90110000000002452c00014697100000e78060169308d00573000000011106ec22e826e44ae02a890869833589016385a5021796010003368629898db3b4c502998013048503086097900000e780001dfd1413040405e5f80335890001cd03350900e2604264a264026905611733000067006373e2604264a2640269056182800c6591c50861173300006700c3718280797106f422f026ec4ae84ee4aa8508612dc903b9050183b98500630b09060144aa840de426846387090003340422fd19e39d09fe814419a80334052151c883598521850497300000e780e06c8355a4212285e3f3b9fe850991cc8e09a29903b50922fd1491c403350522fd14edfc11c8814911a022857d1981442a84e31309fa39a8a2700274e2644269a269456182806387090003350522fd19e39d09fe8335052199c92e8497300000e780c066833504212285e5f911a02a842285a2700274e2644269a2694561173300006700a36497300000e780206417d5ffff1305c5209305b00297800000e78020240000097186fea2faa6f6caf2ceeed2ead6e6dae25efe62fa66f66af26eee2a8a0061ae8a55c883348a008811a2852686d68697100000e780e0ef0e75630605402e7b03b50a0083b50a014e7cee7d2af8aee003b58a0083b50a0203b68a0283bb8a012afc2ef032f463090b080359ab212d45138d0a026376a90c13851d006362a90213060003b385cd02da953305c5025a95b306b9413386c60297800100e78080ec03b50a0193050003b385bd02da9588e903b50a0088e103b58a0088e523bc750103350d0088f103358d001b04190088f5231d8b20a5a603b50a0183b50a00aae02ef803b58a0083b50a0203b68a0283bb8a012afc2ef032f497000000e78000528355a5212d4663ffc5381b861500231dc520130600038666b385c5024276aa9594e9e27690e10276227794e523bc750190f198f52330aa0023340a00054511a622e405491545914c26e863eead006389ad000149994c63979d01814d954c21a0ee8c11a0e51d97000000e780204b8359ab212a8493c4fcffce94231d952013050003b385ac02da9588111306000397800100e7804098314563f6a42c13851c00b385a9406397953013060003b305c502da953386c402228597800100e780a095231d9b2108198c111306000397800100e7806094da8463130900a28452ec03d9a42113851d006362a90213060003b385cd02a6953305c5022695b306b9413386c60297800100e780e0d503b50a0193050003130a0003b385bd02a69588e903b50a0088e103b58a0088e523bc750103350d0088f103358d00052988f5239d242188080c191306000397800100e780a08c03350b216303051481449549a28a835c8b212a8b08018c081306000397800100e780608a631b9c1e835dab212d4563e6ad1a0549114d63ee3c01668d638b3c01014919456395ac00814c154d19a0e51c194d97000000e780603a8359ab212a849344fdffce94231d9520b3054d03da9588111306000397800100e780c084314563faa418930b1d0033857941631e951813050003b385ab02da95130a00033386a402228597800100e780e081231dab2108198c111306000397800100e780a0808359a42113851900b14563f4b9163386ad416316a616050c8e0bda9b93850b22930404220e06268597700100e780a07d014593153500a6958c6133363501239ca5203295b3b6a90093c61600758e23b8852065f288080c191306000397700100e780607a5a856313090022851001e685d68697000000e780a01b03350b21a28ae2849549e31505ec11a0014c97000000e780c02aaa840355a5218145226623b0c42213890422139635004a961062b3b6a500231cb620b6953337b50013471700f98e23389620e5f2c26513851500626a23309a002334aa00639a850d83d9a4212945636c350d1b851900239da420130500033385a90226958c081306000397700100e78040708509139539004a9500e123389420231c342111a810015a85e685d68697000000e780a010626a03350a0105052338aa00f6705674b6741679f669566ab66a166bf27b527cb27c127df26d19618280ad45268531a817d5ffff130535f19305500315a017d5ffff1305d5ed19a8b14597800000e7808065000017d5ffff130575ec9305800297800000e780e0d9000017d5ffff130525d193050002edb717d5ffff130535eaf1bf17d5ffff130585e493050003c9bf17d5ffff1305c5cee9bf83b605219dc683d78521130816009dc71387f7ff93173700b69783b707222330050014e52338050118ed1cf110f50cf92da00ce510e989450ce1828003d7a62119cf03b7862285471ce114e523380501233c05000cf110f518f910fd828097800000e78020ed00001d7186eca2e8a6e4cae04efc52f856f45af05eec62e866e42a84835aa5213689b2892e8a93841500338bba4063e09a0213060003b305ca02a2953385c40222953306cb0297800100e780009e938b1a00130500033305aa02229513060003ce8597700100e780605793892a00130c042213052a00939c3400637c3501b3059c010e05629513163b0097800100e780c099669c23302c01231d742163f434030e0a229a13058a22b305504109461461239c9620850423b88620b38695002105e397c6fee6604664a6640669e279427aa27a027be26b426ca26c25618280411106e413050022c14597300000e780a0ff01c923380520231d0520a260410182801305002297300000e780e0ff0000411106e413050028c14597300000e780a0fc01c923380520231d0520a260410182801305002897300000e780e0fc0000757106e522e1a6fccaf8cef4d2f0d6ecdae8dee4e2e066fc6af8aa8a0075035ca421330bbc002d45636b65112e8983bb8a0183d4ab2163ebb410338a2441239d4b21231d6421130d00033305a90322953306ac03a28597800100e7802089930c1a00338594419305f9ff6318b50eb385ac03de95b309a50322854e8697700100e780e04103b50a0183b40a00330aaa035e9a3305a503aa940a8513060003a68597700100e780a03f130600032685d28597800100e7808083330534018a851306000397700100e780803d83b50a0203b50a03b9c541c9930404220e093385240113163c002106a68597800100e78000808e0ce69b93850b2226854a8697700100e780e0390145050b8c601306150023b88520239ca520a1043285e317cbfe11a031e1aa600a64e6744679a679067ae66a466ba66b066ce27c427d4961828017d5ffff130575c1930530031da017d5ffff1305c5c39305700221a817d5ffff130535b829a017d5ffff1305b5c49305800297800000e78000a50000357106ed22e926e54ae1cefcd2f8d6f4daf0deece2e8e6e4eae06efc2a89033b8501035cab212e8de2952d456363b5148339890203d5a9216364a515b30ca541231dbb20239d9921930bfdff930d00030335090103340900338abb03ae84b38a49013305b5032a940a8513060003a28597700100e780002b130600032285d685a68a97700100e780c06e3305bc035a958a851306000397700100e780a02893041c0033859a406392ab0e3385b4035a95ce85528697700100e780c026b305bd03ce953386bc034e8597700100e780606a8335090203350903adcd4dcd13840922139534005a951305052213193d00a2854a8697700100e780e022b305240113963c002106228597700100e780806663705c030e0c5a9c13058c220c61239c9520850423b865217d1d2105e3180dfe7d556382ac020145938b1c000c601306150023b83521239ca52021043285e397cbfe11a029e1ea604a64aa640a69e679467aa67a067be66b466ca66c066de27d0d61828017d5ffff1305b5ae930520030da017d5ffff1305f5b011a817d5ffff1305959d29a017d5ffff130515aa9305800297800000e780608a0000557186e5a2e126fd4af94ef552f156ed5ae95ee562e1e6fceaf8eef483bd850103dcad21628701c698750357a7216367d71632ec36f02af483ba850283dcaa21130b1c0033069b012d456360c516806188652ae488712ae883bb05010359a42132e0239dcd20130a0003b3844b03a294081813060003a68597700100e780e00f93891b009385040313c5fbff330d250133064d03268597700100e780e05233054c036e950c181306000397700100e780c00c33054b036e9533864c03d68597700100e780800b93050422139539002e9593943b00a695c10513163d0097700100e780804e63f02903a294138584220c611386190023b88520239c35212105b289e317c9fe0315a4217d358545231da420226563f3a50413153b006e951305052293850a2213963c00210697700100e780c00402656372ac02850c0e0c6e9c13058c22da851061231cb62085052338b621fd1c2105e3980cfe626513341500568597300000e78080b27d143375640182752e95a27523b0b501426690e588e9ae600e64ea744a79aa790a7aea6a4a6baa6b0a6ce67c467da67d6961828017d5ffff130515979305100939a017d5ffff1305459f9305a00297700000e780606e0000717106f522f126ed4ae94ee552e1d6fcdaf8def4e2f0e6eceae8eee4033a850183398502035baa2183dba92113041b0033067401ad4563ebc512833c05000c652ee4833d050103ddac2132e0231dca2013090003b38a2d03e69a080813060003d68597700100e78040f593841d0093850a0313c5fdff330ca50133062c03568597700100e780403833052b0352950c081306000397700100e78020f233052403529533862b03ce8597700100e780e0f093850c22139534002e95939a3d00d695c10513163c0097700100e780e03363f0a403e69a13858a220c611386140023b89521239c95202105b284e317cdfe0395ac217d358545239dac20a26463f29504131534005295130505229385092213963b00210697700100e78020ea02656371ab02850b0e0b529b13058b220c61239c8520050423b84521fd1b2105e3980bfe4e8597300000e78060986685a685aa700a74ea644a69aa690a6ae67a467ba67b067ce66c466da66d4d61828017d5ffff130525879305a00297700000e78040560000457186e7a2e326ff4afb4ef752f356ef5aeb5ee762e3e6feeafaeef6ae8483bb050003ba05013289aa8983daab21130b000333046a035e940a8513060003a28597700100e78040df930504031345faff569533066503228597700100e780a022fd3a13950a03239d5b2183ba8400419195456372b51a2819de85568697f0ffffe780a0776a7505cd85456317b5068001080113068003a28597700100e780c0d96a65aa750355a52183d5a5212e950505b1456376b50408180c01014605a88001a80013068003a28597700100e780c0d60675c6750355a52183d5a5212e950505b145637fb5020818ac000546d28697000000e78000bd89a80e65ae6599a0081a13068003a28597700100e780e0d2081a854597000000e78020a03665d66515a0050a081a13068003a28597700100e780a0d0081a854597000000e7804086766596752af82efcd2e0c27be27a03b60b21066a71c293841a00130b010c914d314c954c054d0354a62163e78d0a2819b285268697f0ffffe78040686a750dcd6318a509a81913068003da8597700100e780a0ca526592750355a52183d5a5212e950505636c8503b3858c40a81997000000e780809691a8a81913068003da8597700100e78060c7526592750355a52183d5a5212e95050563728503081a13068003da8597700100e78020c5081a97000000e78020c92a86ae8409a8b3858c40a81997f0ffffe780a079014629fe29a001e405452300a9008a85130600034e8597700100e78060c123b8790323bc590323b04905be601e64fa745a79ba791a7afa6a5a6bba6b1a6cf67c567db67d796182801d7186eca2e8a6e4cae04efc52f856f45af05eec62e866e46ae0b289ae8a2a89938c0601130a0003854b130bf00f03dcaa21b3044c037d54568595cc130d050341055146e68597700100e78060fc932505003335a000b305b040c98d938404fd05046a85e38b75fd13f5f50f631e65016396090089a06284638f09020e045694833a0422fd1965b701452334590123383901233c89002330a900e6604664a6640669e279427aa27a027be26b426ca26c026d256182802334590123380900233c89000545c9bf130101812334117e2330817e233c917c2338217d2334317d2330417d233c517b2338617b2334717b2330817b233c91792338a1792334b1796d71178601001306e6260ce208e61305014997600000e7802060033501497dc98335014a2d466364b6006f10e002138645ff8d4663e4c6006f1040020346d5008346c5000347e5008347f5002206558e4207e207d98f83461500034705008344250003043500a206d98ec2046204458c03388149c18e91445d8e638c960283465500834745008344650003047500a206dd8ec2046204458cc18e8d47e3f5d716f19ac1476397f60063f4c50432856f00507c938605ff8d4763e4d7006f00b07a83461501834705018344250103043501a206dd8ec2046204458c558c931604029b0706008192e362f478e3e3d578b685918d9146e3e7d576f1159306000263fad502154499446306080097200000e780e04e39a08334014a0334814913d58400220593f5f40f4d8d23388148233ca148cda22a968345c6008346b6008347d6008344e600a205d58dc207e204c58fdd8d834606018347f6008344160103442601a206dd8ec2046204458cc18e821633e4b60083454601834636018347560183446601a205d58dc207e204c58f83468601b3e8b7008347760183449601a2060307a600b3e2f600c2048347a6012303e1340307960083458600e207c58f2207d98d2312b13483455600034746008344660083067600a205d98dc204e206c58ed58d2320b13483053602b3e65700821633e91601230cb1388345c6018346b6010347d6018347e601a205d58d4207e207834606025d8fd98d0347f601a2068347160203462602d98e93548900c20762065d8e558e0216d18d2338b1386306080097200000e780a03b0305613483154134032601342303a12e2312b12e2320c12e1305712f0c0f254697700100e7800088135584032307a12e13550403a306a12e135584022306a12e13550402a305a12e135584012305a12e13550401a304a12e135584002304a12ea303812e13d50403230ba12e13d58402a30aa12e13d50402230aa12e13d58401a309a12e13d504012309a12e13d58400a308a12e2308912ea307212f8544e21493851400054597700000e78020801549114409e993852400054597600000e780e07e29cd23382149233c81481305014997f00000e780e0d1aa8413958403619551618330817e0334017e8334817d0339017d8339817c033a017c833a817b033b017b833b817a033c017a833c8179033d0179833d81781301017f82800545621593051500014597600000e780207845c51305014997600000e780a029833d0149638c0d30833c81490336014a13050149ee8597f00000e78080cb13050002814597800000e780c0ab2a8c2e89930501491306000297600100e780c0729305000205460544628597000100e780c0e31375f50f6300052e130501491306004093040040814597600100e780e0622338913805659b08a5811317840305070c0f130501490146814681470148730000006304052ac94429a32334014a2330014a233c014823380148130500022330a13405659b08e5808c061305014989440146814601478147014873000000630295262a840545630ca4241149e31604ea03340134130500020949e36f85e8032501498315414903066149014d2320a1262312b1262303c1260345814983457149034691498346a14922054d8d4206e206558e518d8345c1490346b1498346d1490347e149a205d18dc2066207d98ed58d8215b3eaa5000345014a8345f1490346114a8346214a22054d8d4206e206558e518d8345414a0346314a8346514a0347614aa205d18dc2066207d98ed58d8215b3eba5000345814a8345714a0346914a8346a14a22054d8d4206e206558e518d8345c14a0346b14a8346d14a0347e14aa205d18dc2066207d98e0346f14ad58d82154d8d2300c132233ca130930d1149130c814a1309713a130b11499309814a130a1139fd5c130501490946ea8597600000e78020ec03450149631f053203856d0083855d0003c64d00230ba138a205d18d231ab13803c51d0083c50d0003c62d0083863d0022054d8d4206e206558e518d0334814983158c0003360c008334014a2328a1382314b1342330c1348c0629464a8597600100e780005113558403230fa13813550403a30ea13813558402230ea13813550402a30da13813558401230da13813550401a30ca13813558400230ca138a30b813813d584032303a13a13d50403a302a13a13d584022302a13a13d50402a301a13a13d584012301a13a13d50401a300a13a13d584002300a13aa30f91388c141d465a8597600100e780a048233c51492330714b2c0e25464e8597600100e78040470345013901cd130600025285da8597700100e78060880125630b0512630e9d41050df1b5033581498335014a97f00000e780609685b9014911a0054991b98144ada4833a01391305104063e7aa068545054a568597700000e7804079aa892e84930501491306004097600100e780404093840ac0138509402338913885659b88a58113178a0305070c0f1306004081468147014873000000833501393335a000b3b5b4004d8d31c9e30b04ce4e8597200000e78000ede5b15685814597700000e780c072aa892e8493050149568697600100e780e039914463f19a0222f54545c54b814597700000e78040702a842e8b17b5ffff9305a55899a003c5190083c5090003c6290083c6390022054d8d4206e206558eb364a60022f563989a12a14463f49a1a4545c54b814597700000e780e06b2a842e8b17b5ffff930545544546228597600100e780a032054d1da21305014997600000e780c0a283340149edc0033a81490339014a1305014d13060004814597600100e780c022130541499309014c1306c002814597600100e780602117b5ffff9305f57341464e8597600100e780002d370501011b0505022328a14823340160080f9305014997400000e7804031080fa6854a8697600100e780800e2338a149080f93050149214697600100e780400d233c0134233801342334013423300134130501490c0f1306800f97600100e780e026130501498c061306000297600100e780600b88068c151306000297600100e780406701257dc963070a00268597200000e780c0d41544154989bc033981490334014aa1b44545c54b814597700000e78080592a842e8b17b5ffff9305e5414546228597600100e7804020014d2328a149232a4149233c91482330514b2334814a2338614b233c714b1305014997600000e780608bc9442a7511c54e8597200000e780c0cd63070900628597200000e780e0cce3870c9e6e8597200000e78000ccc5b203c5590083c5490003c6690083c6790022054d8d4206e206558eb364a60013b5840093f53400b335b0004d8d15cd45454544814597700000e780c04eaa84ae8a17b5ffff930525374546268597600100e78080150d4d91bfe30e0a9c268597200000e78080c5f9b263f09a024545c54b814597700000e780e04a2a842e8b17b5ffff93054533c5bb13d524009305f5ff0d4563f0a5044545c54bae8a814597700000e78020482a842e8b17b5ffff930585304546228597600100e780e00e114d8d44e5b517b5ffff1305252b930510026da02ef16398a50a114611444e85d685a68697500000e780e01b13f63500f199b306b5002338a148233cb1482330d14a2334c14a2338814a080f9305014997500000e78000f2080fd68597500000e780801a033401398334013a23388148233c914809452330a14a1305014997500000e780c02b3dc545454544814597700000e780403daa84ae8a17b5ffff9305a5254546268597600100e78000040d4d69aa17b5ffff1305652ef14597600000e780007500004545c54b814597700000e78060392a842e8b17b5ffff9305c5214546228597600100e78020008d44114d8a7aedbbe38504060545e385a406106014644e85d68597500000e780c00d85c12a86ae8613050149b285368697500000e7802012032d014915456314ad100945e38da402106414684e85d68597500000e780600a85c12a86ae8613050149b285368697500000e780c00e032d014915456319ad0c0d45e388a4001068146c4e85d68597500000e780000785c12a86ae8613050149b285368697500000e780600b032d01491545631ead080335813911c5228597200000e78060a593858aff0d456379b54a93854aff6375b54a03c5990083c5890003c6a90083c6b90022054d8d4206e206558eb366a60003c5d90083c5c90003c6e90003c7f90022054d8d42066207598e3367a60013050149ce85568697500000e78060f7833b014a638a0b04833401495e85814597700000e780a0242a842e8aa6855e8697600100e780e0eb0da8032a414983348149833a014a0334814a033b014b833b814b03358139e30f05c80335013997200000e780209a79b101440335814919c50335014997200000e780c098a944e30004ca0d45636475016f10b0010345140083450400034624008306340022054d8d4206e206558e518d85456314b50a13050149a2855e8697500000e7802019033b01498334014a2685814597700000e780001a2a8dae8bda85268697600100e78040e199e06f10607c034b0d0063870b006a8597200000e780e0900335814919c50335014997200000e780c08f63070a00228597200000e780e08e0545054a6303ab000d4a62151306150013050149814597500000e780a070034501491dc1033581498335014a97e00000e780e02caa84f9b6e3060abc228597200000e780808a7dbe031561498315414903562149834611492312a10ec205d18d033481490335814a0356014b8334014aaed1aae9231cc10c6389062e0315410e8e55231aa10a2ed91305610c8c09294697600100e78040d413550403231ea10a13550402231da10a13550401231ca10a231b810a13d504032312a10c13d504022311a10c13d504012310a10c231f910a130501490c19054697000100e780c0a0033401496305042883048149930591491305110f3d4697600100e780e0cda2f52308910e0802ac1197200000e78060c25265930500026304b5006f102069126583451500034605008346250003473500a205d18dc2066207d98ed58d034655008346450003476500834775002206558e4207e2075d8f598e0216d18d2eee83459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2ef283451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2ef683459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5010345f5012206558e42076205598d518d02154d8d2afa130501492c0a528697f00000e780206b03340149630404148304814993059149130511143d4697600100e78060b922fe2300911463070b120545c944631dab4c13050002814597700000e78020efaa842e8b2c0a1306000297600100e78040b6930500020546054a268597f00000e7804027aa8a63070b00268597100000e780406513f5fa0f930450046316454913050002814597700000e78040eaaa842e8b2c0a1306000297600100e78060b1930500020946268597f00000e7808022aa8a63070b00268597100000e780806013f5fa0f854593046004631fb542228597700000e7806006326511c5126597100000e780205e2e7597700000e780e0042a7511c54e8597100000e780a05c63070900628597100000e780c05b63870c006e8597100000e780e05a81446ff0cfac314521a81145b28509a8114539a0114511a03285b68511a0368597700000e780e0a30000b94461b88344814949b883448149c1a6880a2c1a97100000e780607b080f2c1a97100000e780a06f130501492c1a97100000e7804074033401390336013a833401490337014aa812a285a68697e00000e78020060335814911c5268597100000e78000520335813911c5228597100000e7800051080f2c1a97100000e780205f130501492c1a97100000e780c063033401390336013a833401490337014a2803a285a68697e00000e780a0000335814911c5268597100000e780804c0335813911c5228597100000e780804b28132c1a97100000e7802075080f2c1a97100000e780e04d130501492c1a97100000e7808052033401390336013a833401490337014a8803a285a68697e00000e78060fa0335814911c5268597100000e78040460335813911c5228597100000e780404513050149ce85568697500000e78080f08334014a95c0033b01492685814597700000e78080c9aa8bae8ada85268697600100e780c09011a0814b0335814919c50335014997100000e780804063810b1613050149de85268697500000e780c0c3033b01498334014a2685814597700000e780a0c42a842e8dda85268697600100e780e08b23388138233ca1392330913a88060c0f97700000e78040500335814919c50335014997100000e780603a63870a005e8597100000e7808039033501348335813403360135aaf3aef7b2fba8120c191306000297600100e780c0c801259304600263140518130501490c19054697f00000e780a0550334014961c48304814993059149130511203d4697600100e780e082a2ff23009120130501490c19094697f00000e780805203350149aae845c18304814993059149130591213d4697500100e780a07f46652338a120230c9120a81b97100000e780605f9374f50f080c97100000e780805e1375f50f6393a40e080fac1b97100000e780e071130501490c0c97100000e78000710336013a0335014a6311a604833501490335013997600100e78020bc9334150035a0cd44d9a00145814501bb0545854529b30945894511b38344814955a00d458d45e5b98344814979a081440335814919c50335014997100000e780a0260335813919c50335013997100000e7808025a1cc13050002814597700000e78020ab2a8bae8b2c031306000297500100e78040721305014913060002da8597e00000e78020fb0345014959c18344114963870b005a8597100000e780c020466597700000e78080c701a8466597700000e780c0c693047002228597700000e780e0c51e7597700000e78040c55a7511c53a7597100000e780001d766511c5566597100000e780201c7274228597700000e780c0c2326511c5126597100000e780801a2e7597700000e78040c16ff04fcb03358149aae063870b005a8597100000e7806018280e8c1397100000e78040742330012e2338012e280e97100000e7800066aae46308051e814488062c0e268697100000e780006d130501498c0697100000e780405e0335014ad1456304b5006f1060032330014a0335014983451501034605018346250103073501a205d18dc2066207d98ed58d2320b13a83451500034605008346250003473500a205d18dc2066207d98ed58d034655008346450003476500834775002206558e4207e2075d8f598e0216d18d2338b13883459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f83368149598e0216d18d233cb13889c697100000e78000080c0f51461305014a97500100e780e055080f8c0697100000e780403b8335013a4145e39aa5740335013903448500834b9500834aa500034bb5008345c500aef0034ad500034de5008345f500aeec834505002ee983451500aef483452500aefc83453500aef8834545002ef1834555002ee5834565002eed833581390346750032e189c597100000e78040ff8504a20b33e58b00c20a620bb3655b014d8d220a8675b365ba00420d666662063366a601d18d82154d8da675a2054a66d18d66764206c676e206558ed18d2a6622068a76558eea66c2060a676207d98e558e0216d18d2338b148233ca14888159305014997e0ffffe78040960335013497700000e780209f2665e31d95e08335012f0336812e8336012e03358131233cb1222338c1222334d12297700000e780809c03358120833501207e762338a12e2334b12e2330c12e130501498c1597100000e780e0270335014a93050002e31eb5620335014983459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18d2334b13a83451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2330b13a83459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d233cb13883451500034605008346250003473500a205d18dc2066207d98ed58d034655008346450003476500834775002206558e4207e2075d8f83368149598e0216d18d2338b13889c697100000e78000e10335813a8335013a03368139833601392334a14a2330b14a233cc1482338d14888068c1397100000e780c03f080f866597000100e780c09928140c0f13060149940697000100e780e09f058901e90335012e97700000e780c08221a8ae840335012e13f4f50f97700000e7808081e3160442167593050002e310b54cd66703c5970183c5870103c6a70183c6b70122054d8d4206e206558e518d83c5d70103c6c70183c6e70103c7f701a205d18dc2066207d98ed58d82154d8d2334a14a03c5170183c5070103c6270183c6370122054d8d4206e206558e518d83c5570103c6470183c6670103c77701a205d18dc2066207d98ed58d82154d8d2330a14a03c5970083c5870003c6a70083c6b70022054d8d4206e206558e518d83c5d70003c6c70083c6e70003c7f700a205d18dc2066207d98ed58d82154d8d233ca14803c5170083c5070003c6270083c6370022054d8d4206e206558e518d83c5570003c6470083c667003ee403c77700a205d18dc2066207d98ed58d82154d8d2338a148080f9305014997e00000e780404403340139e30c04000335013a83358139130600053306c5022296233081242334b12432e8233cc124e30f05000665930525002eec33b5a5002af0130504052ae1080f13068003a28597500100e7800012087c2aed6307057c03459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8d233ca1260345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8d2338a12603459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8d2334a1260345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8d2330a1266a652330a12828642c0588e5286088e1080597100000e78080eb8275e390051ce2656366b56a130501498c1497e00000e780c0b90335014a2ae56300056a1306814a086a0c6610622330a12c233cb12a2338c12a2a65233ca12808150ce510e188062c0d97100000e78080eb130501498c0697100000e78000e08335014a4145e390a51a03350149034d8500834a95008344a500034ab5008345c5002efc0344d500034be500834bf50083450500aefc83451500aee483452500aef083453500aeec834545002ef183455500aef8834565002ee98335814903467500b2f489c597100000e78020a4a20a33e5aa01c204620ab3659a004d8d2204e275c18d420be20b33e66b01d18d821533eaa50026652205e6754d8d8675c20566666206d18d4d8dc675a2050a76d18d4a664206a676e206558ed18d8215b3e4a500880697100000e78020ce1374f50f880697100000e780e0d733e644018335013493461400558d3364a6002e8597600000e7800043631b04561c1f03c5170183c5070103c627018386370122054d8d4206e206558e518d232ca12c03c5970083c5870003c6a70083c6b70022054d8d4206e206558e518d83c5d70003c6c70083c6e70003c7f700a205d18dc2066207d98ed58d82154d8d2338a12c03c5170083c5070003c6270083c6370022054d8d4206e206558e518d83c5570003c6470083c6670003c77700a205d18dc2066207d98ed58d8215033481224d8d2334a12c833a812333358000033a0123b305a040b3f555012338a148233c01482330814a2334414b2338a14a233c014a2330814c2334414d2338b14c1305014997700000e780a0c269c9aa84130d0501a8055146ea8597500100e780c01c012571fd03250d01906494608c1d88c903350d0088e103358d0088e536e92330d12e32f12334c12e41cc280e9415a285528697e0ffffe78060180335813149e1033501320336813283350133a30f0132630b06368e052e95033505229305f6ff89c90356a5210e06329503350522fd15edf98355a521fd15233ca136233001382334b13813050149ac1e1306f13397e0ffffe780a0ed8806930501491306000397500100e780c0cf0335014c8336014d8355a52163f9b6322a86a9a602e902f1130501490c0597100000e78080b38335014a4145639ca56c03350149834b850003449500034ba500834ab5008345c5002ef4034ad5008344e500034df50083450500aef4834515002ef883452500aee4834535002efc83454500aefc83455500aef083456500aef88335814903467500b2ec89c597000000e780a077220433657401420be20ab3e56a014d8d220aa275b365ba00c204620d33669d00d18d821533e4a50042752205a6754d8da665c20562766206d18d4d8d8675a2056676d18d46764206e666e206558ed18d8215b3e4a500080597100000e78080a11375f50f85456315b502ca65338595003336b5008a76b3858600b2956385d5000a7633b6c500631f065c014a014da1a84a658a7563e385002685ca652e8a63e39500268a8a75638385002a8a0a752a8d63638500228d4a66333596008a76b38586403385a540058e6306d5008a75b3b5a50021a0ca65b3b5c5009386f5ffb3f5a60033f5c600181f104b146718639307014a90cb94e798e3233cb1482338a14828149305014997d0ffffe78080043365aa01630c0514ba757a768806b405980397f00000e78040aa130501498c06054697e00000e78040a7833b014a63800b48033481491306814a08620c66106a833401492330a12e2334b12e2338c12e10070ce608e2233c7137130501498c06094697e00000e78040a3033b014a63030b44033581499305814a906194659869833501492330c12e2334d12e2338e12e181614e710e3269ab3369a003306a4013696233c613163048600b3368600639e0648b345ba00318d4d8d63100540a81e97100000e780208a1374f50f280e97100000e78040891375f50f9304f0076310a43e8815ac1e97100000e780e08c130501492c0e97100000e780008c0336012f0335014a631da600833501490335012e97500100e780a0e61334150011a001440335814919c50335014997000000e780a0530335812e19c50335012e97000000e7808052630d04365a8597600000e78000f95e8597600000e78060f82a6597600000e780c0f76a6597600000e78020f70a652a84c265e317b58a55a82330a134233401342338b134130501498c061306f13397e0ffffe780c0b825a88335814c0336052111ca835685210357a62185053285e3f7e6fe11a0ae86130500033385a60232958c061306000397500100e78080980345f1339385faff233cb122e30c05c8630b0a3c033504222334a1229305faff2338b12223380520228597000000e78080468db983448139f5a40a640da00a652338a12493041004e1a4834401490a652338a12475ac9304b0035da4426423388124880497d0ffffe78080ca880397e00000e780a04a93751500639505208335812203368123b336b00003370123b307d0407d8e2338d148233c01482330b14a2334e14a2338d14a233c014a2330b14c2334e14c2338c14c233c01301b550501233401321dcd931515002e957d15233ca14c1305014997600000e780a07115c1aa85080f1306000397500100e7808089280e0c0f97d0ffffe780a0d70335814d71f5080f0c0c97000000e780c06d0335013a93050002631fb52a0335013983459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18d233cb13483451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2338b13483459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2334b13483451500034605008346250003473500a205d18dc2066207d98ed58d034655008346450003476500834775002206558e4207e2075d8f83368139598e0216d18d2330b13489c697000000e780e026033581358335013503368134833601342334a13a2330b13a233cc1382338d13888158c1397100000e780e08e8806866597f00000e780a0df280e8c06100f941597f00000e780e0e5058911e9280e97d0ffffe78060b029a89b54850039a0ae84280e97d0ffffe78020af13f5f40f49e5281497d0ffffe78020ae466597600000e78000c61e7597600000e78060c55a7511c53a7597000000e780201d766511c5226597000000e780401c72746fe09fbc8344014905a08344014901a8930400085a8597600000e780a0c15e8597600000e78000c10a652338a1242a6597600000e78000c06a6597600000e78060bf880497d0ffffe780009f281497d0ffffe780a0a546656fe0bff71145de856fe05fbd17a5ffff130585d29305b0026fe0efe01795ffff130565536fe00fe017a5ffff130585d89795ffff938625569305b002901497500000e78080ee00001795ffff1305a5506fe04fdd1795ffff1305e54f6fe08fdc41456fe0bfb717a5ffff1305a5d49795ffff938645509305b00213060149c1b717a5ffff130505d39795ffff9386a55065b717a5ffff1305e5d19795ffff9386854f59bf17a5ffff1305c5d09795ffff9386654e51b717a5ffff1305c5db6fe0afcb97400000e780e057000017330000670083c41733000067004301797106f422f026ec4ae84ee43284ae892a89328597300000e78040c2aa8405c163e38900a2892685ca854e8697400100e78080544a8597300000e78060fd2685a2700274e2644269a26945618280011106ec22e826e42a8497300000e78000beaa8401c926858145228697400100e780c0432685e2604264a2640561828017030000670023f717030000670023f717030000670023f717030000670083fb97000000e78080010000411106e497500000e780a0db0000411106e497500000e780c0da0000397106fc22f82a840a850d4697600000e78060d202650dc14265a26502662af42ef032ec2c08228597600000e780a0fce27042742161828017a5ffff130585bd9795ffff9386253d9305b002300897500000e78080d30000397106fc22f82a840a85114697600000e780e0cc02650dc14265a26502662af42ef032ec2c08228597600000e78020f7e27042742161828017a5ffff130505b89795ffff9386a5379305b002300897500000e78000ce0000397106fc22f82a840a85154697600000e78060c702650dc14265a26502662af42ef032ec2c08228597600000e780a0f1e27042742161828017a5ffff130585b29795ffff938625329305b002300897500000e78080c80000397106fc22f82a840a85194697600000e780e0c102650dc14265a26502662af42ef032ec2c08228597600000e78020ece27042742161828017a5ffff130505ad9795ffff9386a52c9305b002300897500000e78000c30000397106fc22f82a840a851d4697600000e78060bc02650dc14265a26502662af42ef032ec2c08228597600000e780a0e6e27042742161828017a5ffff130585a79795ffff938625279305b002300897500000e78080bd0000397106fc22f82a840a85214697600000e780e0b602650dc14265a26502662af42ef032ec2c08228597600000e78020e1e27042742161828017a5ffff130505a29795ffff9386a5219305b002300897500000e78000b80000397106fc22f82a840a85354697600000e78060b102650dc14265a26502662af42ef032ec2c08228597600000e780a0dbe27042742161828017a5ffff1305859c9795ffff9386251c9305b002300897500000e78080b20000397106fc22f82a840a85394697600000e780e0ab02650dc14265a26502662af42ef032ec2c08228597600000e78020d6e27042742161828017a5ffff130505979795ffff9386a5169305b002300897500000e78000ad0000397106fcaa852800014697600000e78080a6226519cd6265c26522662af82ef432f0081097600000e78000c9e2702161828017a5ffff1305e5919795ffff938685119305b002101097500000e780e0a70000397106fc22f82a840a85054697600000e78040a102650dc14265a26502662af42ef032ec2c08228597600000e78080cbe27042742161828017a5ffff1305658c9795ffff9386050c9305b002300897500000e78060a20000397106fcaa852800094697600000e780e09b226519cd6265c26522662af82ef432f0081097600000e780e0b6e2702161828017a5ffff130545879795ffff9386e5069305b002101097500000e780409d0000797106f422f02a840a85194697600000e780a096026519c94265a265026608e80ce410e0a27002744561828017a5ffff130585829795ffff938625029305b0021306f10197500000e78060980000397106fc22f82a840a85094697600000e780c09102650dc14265a26502662af42ef032ec2c08228597600000e78000bce2704274216182801795ffff1305e57c9795ffff938685fc9305b002300897500000e780e0920000397106fc22f82a840a85014697600000e780408c02650dc14265a26502662af42ef032ec2c08228597600000e78080b6e2704274216182801795ffff130565779795ffff938605f79305b002300897500000e780608d0000797106f422f026ec0c6911466394c500814491a0006110600865050610e031c21306450022e06360a6040d4532e46371b504f1152ee80a8597500000e78060740a8597600000e7806080aa84228597500000e78000532685a2700274e26445618280000000001795ffff1305456729a01795ffff1305a5669305b00297400000e780006a0000797106f422f02a840a8597500000e780807e026519c94265a265026608e80ce410e0a2700274456182801795ffff1305656a9795ffff938605ea9305b0021306f10197500000e78040800000797106f422f02a840a85014697500000e780a079026519c94265a265026608e80ce410e0a2700274456182801795ffff130585659795ffff938625e59305b0021306f10197400000e780607b00001d7186eca2e82a842818054697500000e780c074627539c12665866562762aec2ee832e408102c0097600000e7806089027529c14275a2750276aae4aee032fc2c18228597600000e780409d2265e66046642561175300006700a3401795ffff1305a55d9795ffff938645dd9305b002101021a81795ffff1305255c9795ffff9386c5db9305b002301897400000e780207200001d7186eca2e82a842818094697500000e780806b627539c12665866562762aec2ee832e408102c0097600000e7802080027529c14275a2750276aae4aee032fc2c18228597600000e78000942265e6604664256117530000670063371795ffff130565549795ffff938605d49305b002101021a81795ffff1305e5529795ffff938685d29305b002301897400000e780e0680000057186efa2eba6e7cae3ae842a899385050828001306800f97400100e78060d99385040408021306000497400100e78040d803b4841739cc038504001b05f5fb1375f50f1335050c9335140493c515004d8d39e52800a68597000000e780400613060008018e88022295814597400100e78040c788020c02228697400100e78040d328008c021306000897000000e780c00c39a02800a68597000000e78040022c001306800f4a8597400100e78060d0fe605e64be641e693d618280011106ec22e826e44ae02e892a84130505041306800b814597400100e780c0c01795ffff930545c713060004228597400100e78040cc13053900a14522868346e5ff0347d5ff8347f5ff83440500a206d98ec207e204c58f0347150083442500dd8e834735000217a214458fc217830445005d8f1c62d98ee214c58ebd8e14e2fd1521062105c5fd0345090068f4e2604264a26402690561828069ce797106f422f026ec4ae84ee452e03284ae842a89687193050008b389a54063f6c9082330090e130a09065295a6854e8697400100e78040070335090493050508033689042330b904133505f81345150032952334a9044a85d28597000000e78000083304344113051008ce94636fa402930900080335090493050508033689042330b904133505f81345150032952334a9044a85a68597000000e7804004130404f893840408e3e789fc0335090e4a9513050506a685228697400100e780c0fe0335090e22952330a90ea2700274e2644269a269026a45618280417186f7a2f3a6efcaebcee7d2e356ff5afb5ef762f366ef6aeb6ee72e892a842801130600082401814597400100e78040a80d0941458345e9ff0346d9ff8346f9ff03470900a205d18dc206620703461900d98e03472900d58d0216834639002217598e03074900c216558ed18d6217d98d8ce07d15a104210955fd280213060004a28597400100e78080af2c603064833204053267b2772a65aae89756010083b42612033884053e972a97a58db98d9754010083b4641193d605028215d58d338e9500b346fe004a652ae193d78601a216dd8e2a973303d700b345b30013d70501c215b3e8e500469eb345de0093d6f50386055267d274ea67bee4175501000335250db3ebd50026973e97318d398d9755010083b5650c135605020215518daa95ad8c8a7636f813d68401a214d18c3386e600330996003345a900935605014215b36cd500338abc0033459a009355f5030605f26672772a769754010083b44408b369b500ba96b296328c32f433c59200358d9754010083b424079357050202155d8daa94258fca752eec935787012217d98fae96b382f60033c5a200935605014215b36dd500ee94a58f13d5f703860792761666ea75aefc175701000337470333eba700b296ae963345e800358d17570100033767029355050202154d8d2a97398e8e67bef0935586012216d18dbe96b383b60033c5a300135605014215518d2a97b98dae6a13d6f5038605d18d56934e933345a300135605020215498eb29433c53401ce69935685012215c98e338569004ee8b30ed50033c6ce00935706014216336df600b3009d0033c6d0006e6f9356f6030606b36fd6007a99fae033032b01b347130193d407028217c58f3e97b34467010e75aaf493d88401a21433e61401b3086500b298b3c7f80093d40701c21733e39700330be3003346cb002e75aaf81357f6030606b364e600aa92ae9233c69201135706020216598e329eb345be004e7913d78501a2154d8fb30559004af03388e5003346c800935206014216b36256003386c201318fee751355f7030607336ea700ae93ae86aeecde9333c5b301935d050202153365b501b30c4501b3cd7c01926793d58d01a21db3e5bd00be933e873efcb38db30033c5ad00935305014215336a750033059a01a98d93d7f5038605dd8db69eae9eb3c76e0093d607028217dd8e3696b18d93d78501a215dd8db387ee01b38eb700b3c6de0093d70601c216b3e3f6003383c300b345b30013d6f5038605b3ecc500e298fe98b3c5120113d605028215d18d2e953346f501935686012216d18e56e4338658013696b18d93d70501c215b3e8f500b382a80033c5d2009355f50306054d8d4e982698b3450a0193d605028215cd8eb690b3c5900093d78501a215cd8fb3050701b38ff500b3c6df0093d40601c21633e89600c290b3c6f00093d7f6038606d58fca9df29db3c6ad0193d406028216d58c338f6401b346cf0113d78601a216558fe676ee96338ae600b3449a0093d50401c214c58d2e9f3347ef009354f7030607d98c8a66b69eaa9eb3c5be0013d705028215d98d33871500398d935685012215c98e467b33856e01b30ed500b3c5be0013d50501c215b3eba500338deb00b346dd0013d5f6038606b3e0a600466c62963e96334576009355050202154d8d2a9fb345ff0093d68501a215d58d266e7296b309b60033c5a900935605014215558d2a9fb345bf0093d6f5038605b3edd5002676b29fa69fb3c51f0193d605028215cd8e3693b345930093d48501a215cd8c8675fe95b3839500b3c6d30093d70601c216d58f3e93b346930093d4f6038606b3e8960062673a9a669ab3460a0193d406028216c58eb692b3c4920193d58401a214c58d4279b3044901b38fb400b3c6df0093d40601c21633ea9600b3045a00a58d93d6f5038605d58db29eae9e33c5ae00935605020215c98eb382660033c5b200935585012215c98d33855e01b30cb500b3c6dc0013d50601c216b3eea600f69233c5b2009355f50306053363b50033063b010696b18f13d5070282175d8d3388a400b345180093d68501a215d58d62962e96318d935605014215b360d50006983345b8009355f50306054d8dba93ee93b3457a0093d605028215cd8eb387a601b3c5b70113d78501a215b3e4e500b385c301338a9500b346da0013d70601c216b3e3e6009e97bd8c93d6f4038604c58ee275ae9fc69fb3c47f0113d704028214458f3a9fb3441f0193d58401a214c58d827bde9fae9f33c7ef00935407014217458f3a9fb345bf0093d4f503860533ec95008665ae9caa9c33c7ec00935407020217458fba973d8d935485012215c98ce669338599012695298f935807014217336b1701b30cfb0033c79c009357f7030607b36df700ca8a4a96b305d60033c7be009357070202175d8fb307ef00bd8e93d48601a216c58e66762e96338dc6003346ed00135706014216b36ee600338efe00b346de0013d7f603860633efe6000676329a629a33471a00935407020217458fba92b3c5820193d48501a215cd8c8a68b3854801338a95003347ea00935707014217336cf700e292b3c7920093d4f7038607b3e097004267ba9f9a9fb3c77f0093d407028217c58f3e98b344680093d68401a214c58e2279ca9fb69fb3c7ff0093d50701c217dd8db3870501bd8e93d4f6038606c58e329536953346d501935406020216458e33085600b346d80093d48601a216c58e3a953695298e935406014216336396001a983346d8009356f6030606b362d600569d6e9d3346ac01935606020216d18eb69733c6b701135786012216598e3387a801b30ac700b3c6da0093d40601c216b3e39600b38df30033c6cd009356f6030606558e5e9a7a9ab3c5450193d605028215cd8eb3889601b3c5e80193d78501a215cd8fc675d295338ab700b346da0093d40601c21633ef9600fa98b3c7f80093d4f7038607c58fa675ae9f869fb3c66f0193d406028216d58cb38ec401b3c61e0093d58601a216d58db3863f01b38fb600b3c49f0093d60401c214c58eb69eb3c5be0093d4f5038605c58da66b5e953307c500b98e93d406028216c58eb69833c6c800935486012216458e66753a953295a98e93d40601c21633ec9600b30c1c0133c6cc009356f6030606336ed600e26833871a013e9733466700935606020216558e3303d601b346f30093d78601a216dd8e866a5697330dd7003346cd00135706014216598e3293b346d30013d7f6038606b3e0e600ca894a9a2e9ab3467a0013d706028216d98e3698b345b80013d78501a215d98dc66433079a00b38ee500b3c6de0093d70601c216dd8e3698b345b80093d7f5038605b3e3f5006279ca9f969fb3c5ef0193d705028215cd8fbe9db3c55d0013d78501a2154d8f226bb305fb01338fe500b347ff0093d50701c217dd8dae9d33c7ed009357f70306075d8fc2673e953a95298e9357060202165d8e32983347e8009357870122175d8f2695b307e5003d8e135506014216b362a60016983345e8001356f5030605518d2ae8469d729d33c5a601135605020215498eb29d33c5cd01935685012215c98e06756a95330dd5003346cd00135706014216b36fe600338ebf013346de009356f6030606d18ede9e869eb3c5d50113d605028215d18db388950133c61800135786012216598e33873e01b30dc700b3c5bd0093d40501c215b3ee9500f698b3c5c80013d6f50386054d8e569f1e9fb3458f0193d405028215cd8c2693b345730013d58501a2154d8db3052f01b383a500b3c4930093d50401c214c58db3846500258d1357f5030605498f6665aa97b697bd8d13d5050282154d8daa98b3c5d80093d68501a215d58d8a66be96b380b60033c5a000935705014215336af500b30b1a0133c5bb009355f50306053363b50026794a9d329d33c5a201935505020215c98db388b40033c5c800135685012215498e467c33058d01330fc500b345bf0093d70501c215cd8fbe98b3c5c80013d6f5038605b3e2c500667dea9dba9db3c5fd0113d605028215d18d2e983346e800135786012216518f33866d01da89b30ce600b3c5bc0093d40501c215c58d2e983347e8009354f7030607b36f9700c27dee934265aa9333c7d301935407020217d98cb38ac40133c7aa00135587012217598d027e33077e00b30ea700b3c49e0013d60401c214d18c33865401318d9356f5030605558da666b690aa90b3c6f00093d706028216dd8eb38a060133c5aa009357850122155d8db3878001aa97bd8e13d70601c21633e8e600c29a33c5aa009356f5030605b363d5006a9f1a9f33c5e501935505020215c98d2e9633456600935685012215c98e06657a95330dd500b345bd0013d70501c21533e3e500330fc300b345df0013d6f5038605d18d4665aa9c969c33c69401935606020216558eb29bb3c65b0013d78601a216558fb3862c013309d7003346c900935406014216336b9600da9b33c6eb001357f6030606598ece9efe9e33c74e01935407020217d98ca69833c7f801935687012217d98e3387be01330cd700b3449c0013d70401c214458fb3041701a58e13d5f6038606c98e2275aa97ae973d8f135507020217598db30f7501b3c5bf0013d78501a215d98df297338ab7003345aa00135705014215b362e500969f33c5bf008e689355f5030605b369b500469d329d33450d019355050202154d8db30e950033c6ce00ca7d135786012216598eb384ad01338dc4003345ad00135705014215498fba9e33c6ce00926c9357f6030606b36bf60066993699334669009357060202165d8eb29ab3c6da0093d78601a216dd8ee667ca97338ed7003346ce00135506014216518daa9a33c6da009356f60306063369d6008a652e9c1e9c33468b01935606020216d18e369f33467f004e68935786012216d18f33060c01338bc700b346db0013d60601c216558eb306e601b58fae7493d5f7038607dd8dd294ae94258f9357070202175d8f330f5701b3c5e50193d78501a215cd8fb385b401338cb70033478701935407014217336a9700529f33c7e701ca679354f703060733639700ea97ce973d8d135705020215598db303d500b3c6790013d78601a216558fb3869701b30cd70033459501935705014215b369f500ce93334577006e779357f50306055d8d72975e97398e9357060202165d8eb29fb3c7fb014e7e93d48701a217c58f7297338de7003346a601135706014216b36ae600d69f33c6f7012a779357f60306065d8e5a974a97b3c5e20093d705028215cd8fbe9eb345d901ee6693d48501a215cd8cb305d700b382b400b3c7570093d60701c217dd8eb69e33c7d401aa679354f7030607d98ce297aa97bd8e13d706028216d98eb69f3345f501135785012215598dc697330cf500b3c6860113d70601c21633e9e6004ae3ca9f3345f501ea761357f5030605b36be500e696b2963345da00135705020215598d330ad501334646018a7e135786012216598ef696b30dd6003345b501935605014215558d2a9a334646019356f6030606336bd600429d269d33c6a901935606020216558e329fb3c6e401ea6493d58601a216d58db3069d00b38cd50033469601935406014216458e329fb3c5e501ae6493d7f5038605b3e9f500a6929a92b3c55a0093d705028215cd8fbe93b34573008e7493d68501a215cd8eb3859200b38ab600b3c7570193d50701c217dd8db3877500bd8e13d7f6038606d98e629e369e3345c501135705020215598db302e501b3c6560013d78601a216d98e269e338cc60133458501135705014215b363e5009e9233c556009356f5030605336fd5007af6ee98de9833451601135605020215518d3303f50033c66b00ee76135786012216598ec696b30bd60033457501935605014215336ed5007293334566002e769356f5030605558d66965a96b18d93d605028215d58db386f5013347db00ca67935487012217d98c3e96338bc400b3c5650113d60501c215b3efc500fe96b58c93d5f4038604b3ecb400d69ece9eb345d90113d605028215d18d2e9a33c64901935486012216d18c33860e01b38ac400b3c5550113d60501c215d18d2e9a33c64401ca741357f6030606598ee294aa94a58d13d705028215d98dae96358d2a679357850122155d8d2697330de500b3c5a50113d70501c215b3eee50076e3b388de0033451501126c9356f50306053369d500e29be69b33c57301935605020215c98eb383460133c57c002a77935785012215c98f3385eb00338aa700b3c6460113d70601c216558fba93b3c677002e6893d7f6038606b3ebf600429b329bb3466e0193d706028216d58fbe9233465600ea75935686012216558eb306bb00330bd600b3c7670113d50701c2175d8daa92334656006a6e9357f6030606b369f600f29afa9a33c65f01935706020216d18f3e9333466f00ee66935486012216d18c3386da002696b18f93d60701c217dd8e3693b3c7640093d4f7038607c58fea95be952d8f935407020217d98ca69233c75700935787012217d98fe295b38ab700b3c4540193d50401c214b3efb400fe92b3c5570093d7f503ee74860533eff5007af6d294ca94258d935505020215c98d2e9333456900ce67135785012215498f3385f400330ca700b3c5850193d70501c21533eaf5005293b34567000e7793d7f5038605cd8f5a975e97b98e93d506028216d58dae98b3c61b018a7413d58601a216558d2697b304e500a58d93d60501c21533e9d500ca9833451501aa659356f5030605558db295ce9533c6be00935606020216558eb293b3c6790013d78601a216d98ec2953388b60033460601135706014216598eb293b3c676002e7793d5f6038606d58d56973e97398e935606020216558eb298b3c6170193d78601a216d58fb306c701b389d70033463601135706014216b36ee60076e3f69833c617014e779357f6030606336bf60062972a9733c6ef00935706020216d18fbe93334575008e6f135685012215518d3306f701330cc500b3c7870113d70701c2175d8fba93334575004a6e9357f5030605b36af500f294ae9433459a009357050202155d8daa92b3c555002a7a13d68501a215d18dd294b38c950033459501135605014215336dc500ea92b3c555006e6693d6f5038605b3ebd50032987a98b345090193d605028215cd8eb3846600b3459f004a7393d78501a215cd8fb30568003389b700b3c6260193d50601c216d58dae94a58f93d6f7038607dd8e4e963696318f9357070202175d8f33085700b3c60601ea6713d58601a216558d3e96b30dc5003347b701135607014217b369c7004e98334505011356f5032e670605336fc5007af662975a973345ed00135605020215518db302950033465b009357860122165d8e5297330be60033456501135705014215336ae500d292334556001356f5030605518de69fd69fb3c5f50113d605028215d18d3387150133c6ea00ea74935786012216d18f33869f00b38fc700b3c5f50193d40501c215b3e895004697b98f93d5f7038607dd8d4a9e5e9eb3c7ce0193d407028217c58fbe93b3c47b0013d68401a214458e7293b30e6600b3c7d70193d40701c217c58fbe933346760092649356f6030606558eee94aa94a58f93d607028217dd8e3383e600334565000e779357850122155d8d2697b30be500b3c6760193d70601c21633eef60072e3729333456500ce669357f50306053369f500da96ae9633c5d900935705020215c98fbe9333c57500ee75935485012215c98c3385b600338ba400b3c7670193d50701c217dd8dae93b3c674008a7a93d7f6038606b3e9f600d69fb29fb346fa0193d706028216dd8e369833460601ae77935486012216458efe97330cf600b3c6860193d40601c216c58e369833460601ce741355f6030606336aa600a69efa9e33c5d801135605020215518daa9233465f002a67935486012216458eba9e330fd6013345e5019357050142155d8daa92334656009357f60306065d8e5e973297b98d93d705028215dd8d2e9833460601ca67935486012216d18c3306f700b38cc400b3c5950113d70501c215b3efe5007e98b3c5040113d7f503ea678605b3eee50076f6da97ca97bd8e93d506028216cd8eb3885600b345190113d78501a2154d8fb3855701330bb700b3c6660193d70601c216b3eaf600d69833471701aa779354f7030607458fe297ce973d8d935405020215458d2a93b3c46900ca7693d58401a214c58dbe96b38bd500334575019356050142153369d5004a9333c56500ea759356f5030605c98efa95d2953345be00935405020215c98ca69333457a008e67135685012215498e3385f500330ca600b3c4840193d50401c214c58db38775003d8eae629354f6030606458e969cba9cb3c5950193d405028215c58db3836500334777004e63935487012217458fb3846c00330d9700b3c5a50113d50501c21533efa500fa9333457700ee6c9355f5030605b369b500669b369b33c56f019355050202154d8daa97bd8e8e7513d78601a216d98eda95338bb60033456501135705014215498f330ef70033c5c601ae769357f5030605336af500de96b29633c5da009357050202155d8d2a9833460601ce7f935786012216d18f3386f601b38bc70033457501935605014215558d2a98b3c50701ee7793d6f5038605b3ead5003e9c769cb345890193d605028215d58dae98b3c41e01926613d68401a214458eb304dc0033099600b3c5250193d40501c215c58dae98334616019354f6030606458eea97b2973d8f935407020217458f3a9833460601935486012216458ee697330cf60033478701935407014217b36e97007698334606011357f6030606aa74598e7ae332f6da94ce94258d135605020215518d3306150133c7c900935787012217d98f33875400b389e70033453501935405014215b36895004696b2ea3d8e1355f6030606b367a6005e93529333c565009355050202154d8daa93b3457a0013d68501a215d18d3306d3003383c50033456500935605014215b362d500969333c575009355f5030605b366b500ca9fd69f3345ff01935505020215c98d2e9e33c5ca01ea74135685012215498e33859f00330fa600b3c5e50193d40501c215cd8c269eb345c6014a6613d5f5038605c98d62963e96b18c13d504028214458daa93b3c77700ae7413d78701a2175d8f26963a9632e6318d135605014215518d2ae31e95aaee398d1356f5032a670605518d2afa4e97369733c5ee00135605020215518d2a9e33c6c601ea669357860122165d8eba96b29636ea358d935605014215558daaf67295aaf2318d1356f5038e760605518d2afe9a96ae9633c5d800135605020215518d2a98b3c505010e6613d78501a215d98d36962e9632ee318d135605014215518daafa4295aae62d8d9355f50306054d8daae23275ca75aa95fa9533c6b200d666135706020216598eb296358d0a779357850122155d8dba95aa952ef2b18d13d60501c215d18daefeb695aeea2d8d9355f5030605c98da8022ef6a1451060833605fc1861358e398e10e0fd1521052104f5f5be701e74fe645e69be691e6afa7a5a7bba7b1a7cfa6c5a6dba6d7d6182801d7186eca2e8a6e4cae02e89aa840a8513060004814597200100e780a0fae8749305000263e9a50aa86855e5e870ac603386a500b46403c7040fb335b600b0e0b695ace419c3fd55acecfd5513061008ace86378c50813060008138404066309c500098e2295814597200100e78080f52685a28597e0ffffe780e04921459305310026861462a38ed5fe13d78600238fe5fe13d70601a38fe5fe13d786012380e50013d70602a380e50013d786022381e50013d70603a381e500e1922382d5007d152106a1055dfdf0748a854a8597200100e78000fce6604664a6640669256182809305000897300000e78020f70000657106e722e3a6feae842a84938505080a851306800f97200100e78080f8a81913060004a68597200100e78080f793850404281a1306000497200100e78060f683b6841789ca0a85ac19301a97200100e78040d439a00a85ac1997200100e78040c98a851306800f228597200100e78040f3ba601a64f67459618280197186fca2f8a6f4caf0ceecd2e8d6e4dae05efc62f866f46af06eec906103bc8500329c636fcc34aa8988699376f50093b616003337a000f98e6380063a814a89466368d5008d462a87850a0581e3ede6fe83cb85013285d68597000000e780a03b6365ac322a8d1305000463f5aa323305ac4133555501814c89456368b5008d452a86850c0581e3edc5fe938d2c0063ea9d316145b3b5ad02639a0530b384ad02ea9463eaa43113893c006a847d19268a630d0902630c0d24233044015285639b0b00130600105285814597200100e78080d80860610408e1c10408e5e3f844fd1775ffff130525f0a5ac4ee0638b0d2e014b13098d0093891c005a85ee8597000000e780a03563030d201d05935435002330490163990b0052858145268697200100e78040d3d29463e24425638669016109050b268ad1b7094963e72d0593098d02330a904105442285ee8597000000e780c0301d05135b350023b0990063990b00268581455a8697200100e780a0ce33856401636195200504b3058a00e109aa84e39325fd11a02685d68597000000e7806028636fac2463860d262a8b938bfdff2a84638b0b161385edff9305f00363eda520854c5a846ae86ee463080d14aa843395ac00331d55013309a401636589186145b38da402c265ae9d3385ab022e9593098500130a0501636f2c0d03b50d000c612300b40013d68503a303c40013d605032303c40013d68502a302c40013d605022302c40013d68501a301c40013d605012301c400a181a300b40093558503a307b400935505032307b40093558502a306b400935505022306b40093558501a305b400935505012305b40093558500a304b4002304a4000c6180e500e15a85d6852686a28697000000e780c022058915ed5a85d6855e86a28697000000e780802183b5090013563500b295838605001d893395ac00c98e2380d50083350a00b29503860500518d2380a5004a846a99e37489f249a82685a26597000000e780c0185a85d6852686a28697000000e780801c83b58d0013563500b295038605001d893395ac00518d2380a50081cc1385f4ffa68b426de31c0dea97200000e780804f0000426da26d63638c0a33058c40826523b0650123b4850188e923bca50123b0b50323b45503e6704674a6740679e669466aa66a066be27b427ca27c027de26d096182801775ffff1305a5c8f14597200000e780402e00001775ffff130565c7f5b71775ffff1305c5c6cdb71775ffff130525c6e1bf1775ffff130585bfada81775ffff1305e5c193054002c9b71775ffff130505c45dbf1775ffff130565baa1a81775ffff1305c5c24db71775ffff130525bc91a01775ffff130585b59305300271b71775ffff1305a5c429a85285d68597000000e780c002637bac001775ffff130585c797000000e780400500001775ffff1305e5b79305100289bf01cd1306000463f0c5027d153355b50005053315b50082801775ffff130585b59305100239a01775ffff1305a5b79305400297200000e7802020000097200000e780403c000063efa5006382a5021345f5ffaa951305000463f2a50205453315b50082801775ffff1305c5b029a01775ffff130525b09305100239a01775ffff130545a99305300297200000e780c01a000063e0a6041307f003636cc7001307000463fde500898e33d5c6003355b50082801775ffff1305e5ae29a01775ffff130545ae9305400297200000e780c01600001775ffff130565b9b545f5b790659461137806fc3698636bd80c98699355660063e3e500ba8594e2094694e6b68763ebc508fd1593d8860393d2060313d3860293d3060213de860193de060113df8600b68736863e879387070463efe7062380c70013578603a383e700135706032383e70013578602a382e700135706022382e70013578601a381e700135706012381e7002182a380c7002384d700a387170123875700a386670023867700a385c7012385d701a384e70190621ce6fd159ce23e86c9f99385070463e7f50214e1233405010ce914ed82801775ffff130565a2f14597200000e780000800001775ffff130525a1f5b71775ffff130585a0cdb7717106f522f126ed4ae94ee552e1d6fcdaf8def4e2f0e6eceae82a841305000497350100138ae5ff6371850417350100930425ff8860631e05348864fd558ce063130512c870cc6cd068d464aae4aee032fc36f80a850c1897000000e780209c054588e413850401c5a803350a04631b053203358a04fd552330ba041ded03350a0883358a0703360a07aae02efc32f80a850c1897000000e78080e705452334aa040265a2654266e2662338aa04233cba042330ca062334da0603398a0663000902033509000c6110650ce20c6510610ce6130b0a04630825032a8991a403390a0603358a056373a902130509046368252983350a042330aa0685052330ba046315092209a823340a0619ac03350a0405052330aa0403350a00631e052803358a00fd552330ba001ded03350a0a83358a0903360a0983368a08aae4aee032fc36f80a850c1897000000e780408d05452334aa0013050a018a851306000397100100e780e07d83398a031305f003636335210545814c3315350163788500850c63840c1c0605e36c85fe83350a0363e3bc00e68503358a020146e146b386dc02aa96138406fdb385bc406389c516630d051c147803b9060061047d16e307d9fe033509008335890088e1033589008335090088e5047017350100130b85e403350b0183358b03934af6ffe69a5686ca8697000000e78000cd93553500a695038605001d89854b3395ab00518d2380a50063f85c11130c000417350100130b65e0138afaff63778a1333954b01b3143501ca9463e72413033d840203350b0183358b035686ca8697000000e780a0c793553500ea95038605001d893395ab00518d2380a500833a840003350b0183358b035286ca8697000000e780c0c493553500d695038605001d893395ab00518d2380a50008600c612380b40013d68503a383c40013d605032383c40013d68502a382c40013d605022382c40013d68501a381c40013d605012381c400a181a380b40093558503a387b400935505032387b40093558502a386b400935505022386b40093558501a385b400935505012385b40093558500a384b4002384a4000c6184e504e12114d28ae3e54cf119a00149528b03350b0005052330ab004a85aa700a74ea644a69aa690a6ae67a467ba67b067ce66c466d4d6182801765ffff1305656b21a81765ffff1305c55e9305300231a01765ffff1305e569f14597200000e78080cf00001765ffff1305a55cf9bf1765ffff13050568cdb797200000e78080e900001775ffff1305d5a19765ffff9386455815a01775ffff1305b5a09765ffff9386255709a81775ffff1305959f9765ffff93860556c1450a8697200000e78080e40000317106fd22f926f54af14eed52e956e55ae1defce2f8e6f4eaf0eeec97350100938ce5c283b50c04639d05382a8903b58c04fd5523b0bc041de917350100130405c148602c7c3078aae4aee032fc28002c1897000000e78060ae054528e42265c2656266827628e82cec30f034f403b50c0583b58c053335a9001345f5ffb335b9006d8d51c517350100130545bc2c75638e052090612300c90093568603a303d900935606032303d90093568602a302d900935606022302d90093568601a301d900935606012301d9002182a300c90013d68503a307c90013d605032307c90013d68502a306c90013d605022306c90013d68501a305c90013d605012305c90013d68500a304c9002304b900906165a203b50c0483b50c00050523b0ac04639b052a03b58c00fd5523b0bc0015ed173501001304c5b148704c6c50685464aae8aee4b2e036fc28002c1897f0ffffe780c04f054508e4130504012c001306000397100100e780804083ba0c03638f0a2283b98c02138afaff13848902854463809a04638b0922033b040003b50c0183b58c032686ca8697000000e780609593553500da9583c505001d8933d5a50005898504610469d5f91463e6440139a263030a108144930a0004268b63e49a00130b000483bb8c0303bc0c0161453385a4024e9513048502054d03b50c0183b58c032686ca8697000000e780808f638e091a833504fe13563500b2950386050093767500b316dd0093c6f6ff758e2380c500937515003306b040833604fe13661600329513563500369603460600937675003356d600058a51e2630b9b1263fe5b1333159500331575016295636e85131061146590e21065146190e691c12a89833d040003b50c0183b58c0385042686ca8697000000e780c08693553500ee95038605001d893315ad001345f5ff718d2380a5006104e3129af4d28405a023302901930585064a862334260123b02501930c050451a8638a090e814461453385a4024e9508610c612300b90013d68503a303c90013d605032303c90013d68502a302c90013d605022302c90013d68501a301c90013d605012301c900a181a300b90093558503a307b900935505032307b90093558502a306b900935505022306b90093558501a305b900935505012305b90093558500a304b9002304a9000c6123b425012330250103b50c00050523b0ac00ea704a74aa740a79ea694a6aaa6a0a6be67b467ca67c067de66d296182801765ffff1305c51e29a01765ffff1305251e9305300231a01765ffff13054529f14597200000e780e08e00001765ffff1305052293051002edb797200000e78040a900001765ffff130595619765ffff9386051809a81765ffff130575609765ffff9386e516c145300097200000e78060a500005d7186e4a2e026fc4af84ef452f056ec83ba050263800a0a2e8a2a898065b35954034e8597000000e780200b83340a002ae02ee402e863e335078145636e54031396350032950d466370560983c6140003c70400a206d98e03c7240083c7340033045441d6944207e2075d8fd98e14e185052105e37a54fd2ee8226502662338b9002334a9002330c900a6600664e2744279a279027ae26a616182800a8581454e8697000000e7806008c2650265e37954f9d9b71765ffff13054523e54597100000e780e07d00001145d68597200000e78040070000011106ec22e826e42a841dc51355c40305ed93351500931434008e0599c4268597d0ffffe780a0b8aa8581e9268597d0ffffe780c0b90000a1452e85a285e2604264a2640561828097d0ffffe780c0b80000411106e497000000e78000037d567e1605066315c500a2604101828011e597d0ffffe78040b600002e8597d0ffffe780e0b400005d7186e4a2e026fcae86b29563f4d5000145a1a82a8408659314150063e39500ae84914563e39500914493d5c40393b51500139634008e0501c914600e0536f0a14636f42af811a002f42800141097200000e7800028a265426599c1e26531a008e004e47d557e150505a6600664e27461618280411106e4054697000000e78060f87d567e1605066315c500a2604101828011e597d0ffffe780a0ab00002e8597d0ffffe78040aa0000797106f422f026ec4ae84ee452e06365d7046366e604aa89b304d7403389d5002685814597200000e780802c2a842e8aca85268697100100e780c0f323b0890023b4490123b89900a2700274e2644269a269026a456182803685ba8519a03a85b28597200000e78080ed000063e8c60063e9d500b385c640329582803285b68511a0368597200000e78060eb0000011106ec22e826e42a8410690865ae846319a6002285b28597000000e78040f210680860931536002e9504e1050610e8e2604264a26405618280397106fc22f826f44af04eec52e856e4114a32892a84637d46032d45ad4a814597200000e7804020aa84ae891765ffff930505042d46268597100100e78000e7054508c0233444012338240104ecb1a803c5150003c6050083c6250083c535002205518dc206e205d58db3e4a500b9c09104638424052d45ad4a814597200000e780801a2a8aae891765ffff930545fe2d46528597100100e78040e12320040004e423382401233c4401233034032334540331a0114a631d4901154508c0e2704274a2740279e269426aa26a216182802d45ad4a814597200000e780e014aa84ae891765ffff9305a5f82d46268597100100e780a0db23200400a9b71061833805011c65210605483e8763ee17019307f7ff10e11ce5637d1801833686ff0c622106e3f3d5fe333517011345150082800545854597200000e780e0d30000797106f422f026ec4ae84ee452e02e89aa8413050002130a0002814597200000e780a00c2a84ae8913060002ca8597100100e780c0d380e023b4340123b84401a2700274e2644269a269026a45618280397106fc22f826f44af0b2841106636996042e892a843285814597200000e780c0072ae02ee402e826ce10100a856c0897200000e780e0ec330699000a85ca8597200000e780e0eb4265a265026608e80ce410e0e2704274a2740279216182801765ffff1305c5e4f14597100000e780603d0000797106f422f026ec4ae84ee452e08d4663f3c604aa899304c6ff138945002685814597200000e78000002a842e8aca85268697100100e78040c723b0890023b4490123b89900a2700274e2644269a269026a456182801145b28597200000e78060c10000011106ec22e826e44ae02a841305000285451309000297c0ffffe780607329c9aa8413060002814597100100e780c0b404e0233424012338240111458545914497c0ffffe780c0701dc5a301050023010500a30005002300050008ec04f004f423080402e2604264a2640269056182801305000211a0114597c0ffffe780406f0000757106e522e1a6fccaf8cef4d2f0d6ecdae8dee4e2e003bb050193040b0163e86415938b140063890b142e8a83ba8502b3895b0163e779152a894e85814597200000e780e0ef2ae42ee802ec0d4597000000e78020ad2af02ef402f899c1814501a8081097000000e78060bbc27502758e052e95c1450ce1c27585052ef822756398a500081097000000e78040b9c275027c13953500629504e19384150026f82275639aa4000810a68597000000e78000b7c274027c1394340033058c00233075014ede900028006c1897200000e780a0cda2797d556384a402930b0104210462850c61930485002ede28006c185e8697200000e78040cb611426857df063870900628597c0ffffe780e05c83350a0013040a0333866501280097200000e780a0c813061a032800a28597200000e780a0c783358a0133865501280097200000e78080c66265c26522662338a9002334b9002330c900aa600a64e6744679a679067ae66a466ba66b066c496182801765ffff130545be11a81765ffff1305a5bd29a01765ffff130505bdf14597100000e780a01500000d476371c7069306c6ff637ad704930686ff0d476375d70403c8550003c7450083c7650083c6750022083367e800c207e206dd8ed98e03c8950083c8850083c2a50083c7b500220833671801c202e207b3e757005d8f17030000670043a61145b68519a01145b28597200000e780c0980000411106e410610e069766ffff93862681369610620286907588711c6e9765ffff938595c33d4635a8907588711c6e9765ffff9385c5c12d462da021052ae01765ffff9307c5bd1765ffff130745be3d463da0907588711c6e9765ffff9385a5ba2146a2604101828721052ae01765ffff9307b5b61765ffff1307e5b61d468a862e85be8597200000e7806086a2604101828082808365050005466345b60099c9054609a809466389c5000d466394c500210521a0610511a041050c6591c5086117c3ffff6700a3408280130101ba233c1144233881442334914423302145233c3143233841432334514323306143233c71412a8b08081306004013040040814597000100e780a07e2338814005659b0895819305014105470808014681468147014873000000aa84094505446384a412638084081144639f0410033a0141130500406379450785450544528597200000e78080beaa892e890c081306004097100100e780a08593020ac0138509402338514085659b88958193050141130600400547094381468147014873000000630c650aaa846308850a1144d5e483340141094463e2920a13054afd1334150035a001444da05285814597200000e780c0b7aa892e890c08528697000100e780007f1305c00201446306aa023d45bd4b814597200000e78040b5aa84ae8a1765ffff9305b59c3d46268597000100e780007c01c823303b0123342b0123384b0189a802c81305c0022aec52f026f456f85efc0d452334ab0023300b00080897000000e78080e6630609024e8597c0ffffe780002939a80144630709004e8597c0ffffe780e02723348b0023389b0023300b008330814503340145833481440339014483398143033a0143833a8142033b0142833b8141130101468280397106fc22f83287ae862a8402f002ec02e802e4130500022af405659b0815822c108d472800894201460148730000006309550285456308b502914515e522751306000289456361a602130514002c001306000297000100e780a06d2300040009a8854511a081450ce408e805452300a400e270427421618280397106fc22f83287ae862a8402f002ec02e802e4130500022af405659b0815822c109547280089420146014873000000630b55028545630cb502914515e922751306000289456365a602130524002c001306000297000100e780006601458545a300b40009a80145a300040029a081450ce408e805452300a400e270427421618280130101ba233c1144233881442334914423302145233c3143233841432334514323306143233c7141b289ae8b2a8408081306004093040040814597000100e780a0522338914005659b08c58293050141080889440146de864e8781470148730000006301950885456300b508914535ed03390141130500406372250b8545054b4a8597200000e780c0922a8aae8a0c081306004097000100e780e059930209c013050a402338514085659b88c58293050141130600408944de864e87814701487300000063019508630e6507114b25ed03350141094b63e8a2062330440123345401b1a8854511a081450ce408e8233004008330814503340145833481440339014483398143033a0143833a8142033b0142833b81411301014682804a85814597200000e780e088aa84ae890c084a8697000100e780205004e0233434012338240145bf014b2334640108e823300400e3810afa528597c0ffffe780e0fe51bf130101b8233c1146233881462334914623302147233c3145233841452334514523306145233c714323388143233491432330a1432a8d28001306004013040040814597000100e780203c2334814005659b08458093058140280009440146814601478147014873000000aa84630f85060545638ea4061144639b0412833b81401305004063777507854505445e8597100000e780007caa892e892c001306004097000100e780204393820bc0138509402334514085659b884580930581401306004009438146014781470148730000006308650caa846304850c1144f1e083348140094463ee920aa1a00544c9a001447da85e85814597100000e7808075aa892e892c005e8697000100e780c03c114a63f04b033145b14c814597100000e7804073aa8a2e8b1755ffff9305f55925aa03c5190083c5090003c6290083c6390022054d8d4206e206558e336aa60063934b03214a63fe4b093145b14c814597100000e780006faa8a2e8b1755ffff9305b555d5a83145b14c814597100000e780406daa8a2e8b1755ffff9305f5533146568597000100e78000348144e1a80144630709004e8597c0ffffe780e0e323348d0023389d0023300d008330814703340147833481460339014683398145033a0145833a8144033b0144833b8143033c0143833c8142033d014213010148828003c5590083c5490003c6690083c6790022054d8d4206e206558e336aa60013358a0093753a00b335b0004d8d15c53145b14a814597100000e780a0622a8aae8b1755ffff930555493146528597000100e78060298d443da063ff4b053145b14c814597100000e780c05faa8a2e8b1755ffff930575463146568597000100e7808026854426c462c652e85eec56f05af466f80d452334ad0023300d00280097000000e7800092e30209f24e8597c0ffffe78080d419bf13542a007d140d456379a4023145b14c814597100000e7806059aa8a2e8b1755ffff930515403146568597000100e78020209144a28b0d4a59bf6316a408114611444e85de85d28697f0ffffe780002e13f63500f199b306b5002ae42ee836ec32f022f4130581402c0097f0ffffe780c00413058140de8597f0ffffe780202d833a81400334814156e422e809452aec280097f0ffffe780e03e29cd3145b14a814597100000e78060502a8aae8b1755ffff930515373146528597000100e78020178d4411aa3145b14c814597100000e780c04daa8a2e8b1755ffff930575343146568597000100e780801491440d4aa28bf1bd6304041005456304a41003b60a0083b68a004e85de8597f0ffffe780e021130a0002639b450709456306a40e03b68a0083b60a014e85de8597f0ffffe780c01f054a639b45070d456309a40c03b60a0183b68a014e85de8597f0ffffe780c01d2a86ae862800b285368697f0ffffe7806022a24415456392a4080335014111c5568597c0ffffe78080bc23303d0123342d0123387d0169b32e8c3145b14c814597100000e7804041aa8a2e8b1755ffff93054524314605a02e8c2945a94c814597100000e780403faa8a2e8b1755ffff9305a5212946568597000100e78000068144e28b03350141e30905de0335814097c0ffffe780a0b5cdb3324c426ae26b827a227bc27cf9bf0145814509a80545854531a00945894519a00d458d4597100000e78040fe00009308d0057d558145014681460147814701487300000001a041112e87aa8602e405659b0875812c000545014681470148730000001335150041018280086101a08280797106f42e8813564500130f7002130710279756ffff938ee62e6363e608130f700213076102171601008338a66239661b03068f05669b03b6479302c0f937e6f5051b0ef60faa86333515032d813b066502b307d600139607034992330676029355160141821376e67fbb855502be95769683471600c615c19103460600a30ff7fef69583c7150083c50500711f230fc7fea300f7002300b7007117e365defa130630066370a60493150503c99105661b06b647b385c502c5811306c0f93b86c502329546154191791f7695034615000345050093061100fa96a380c6002380a6002e85a945637cb5009305ffff130611002e961b0505032300a60005a006059305efff7695034615000345050093061100ae96a380c6002380a60093061100ae96130770020d8f1755ffff9305855d4285014697000000e780e000a27045618280597186f4a2f0a6eccae8cee4d2e056fc5af85ef462f066ec6ae86ee4aa8403654503ba893689328aae8b937c1500b70a110063840c00930ab00293754500ce9c89e5814b8c6085e5a1a08145630e0a005286de86038706008506132707fc134717007d16ba957df6ae9c8c6095c103bd840063ffac01218925ed83c58403054633059d41634cb60af9e1aa8c2e85c9a0807084742285a6855686de86528797000000e7806014054b0dc15a85a6700674e6644669a669066ae27a427ba27b027ce26c426da26d656182809c6c2285ca854e86a6700674e6644669a669066ae27a427ba27b027ce26c426da26d6561828780581305000383c584032ee003bc040283bd840288d8054b238c64036285ee855686de86528797000000e780e00c51f5228a33049d4105047d1451c803b60d02930500036285029665d985bf09466398c50093051500058193dc150011a0814c03bc040203bd84028458130415007d1409c803360d026285a68502966dd9054b2dbf37051100054be389a4f26285ea855686de86528797000000e780e00511fd83368d016285ca854e86829619f5b30990417d5a7d59338529016309450303360d026285a6850296050975d50da083b68d016285ca854e868296e31005ee014b23a844030265238ca402c1bd6689333b9901e1b5797106f422f026ec4ae84ee49b070600370811003a89b6842e84aa896389070114704e85b2858296aa85054591ed81cc1c6c4e85a6854a86a2700274e2644269a269456182870145a2700274e2644269a269456182805d7186e4a2e026fc4af84ef452f056ec5ae85ee483320500146933e7d2003289ae896304072a638706101c6d8146338e29018507370311009308f00d1308000f4e8601a893051600918eae962e866303640efd17adc7630fc60d8305060013f4f50fe3d105fe834516009374f40113f7f50363fa8802834526001a0793f5f503b363b7006367040383453600f614ad909a0393f5f50333e4b300458c630c64089305460055b79305260013946400598c61bf93053600b20433e4930071b7630bc6078305060063d3050493f5f50f1307000e63ede5021307000f63e9e50203471600834726001377f70393f7f70303463600f615ad9132079a075d8f1376f603598ed18d370611006386c50285c263fd2601b385d90083850500130600fc63d7c500814591e539a0e39d26ffce8599c13689ae89638b021803388500930500026372b902814e63060916ca85ce86038606008506132606fc13461600fd15b29efdf581aa13877900619b3386e940b308c90093f678008145630d3701ce87038407008507132404fc934414000506a6957df6014691ce93f788ffba9783840700850793a404fc93c41400fd162696fdf693d638009717010083b787129714010083b28412b714001092048504939804018508b30eb6001da013173e001a97b386c34113763e00b3f45500a181b3f55500a695b3851503c191ae9e2deaddcab6833a839305000c368e63e4b600130e000c9375ce0f139435001a94dddd81451a8745df146393c4f6ff9d8099821067c58efd8eb6959346f6ff9d82046b1982558e7d8e93c6f4ff9d829980c58e046ffd8e3696b29513c6f4ff1d829980458e7d8e13070702b295e31d87fabdb7630803029305000c63e4b3009303000c814593f633008e06106021041347f6ff1d831982598e7d8ee116b295f5f611a0814533f65500a181b3f55500b295b3851503c191ae9e63fc0e01834685030546b305d8416345d60285ce814a25a80c7508719c6dce854a86a6600664e2744279a279027ae26a426ba26b6161828709466398c600138615008581935a160019a0ae8a8145033b0502833b85020459138415007d1409c803b60b025a85a68502966dd9054a81a037051100054a638ca40283b68b015a85ce854a86829605e533095041fd597d5433058900630a350103b60b025a85a6850296050475d511a05684333a54015285a6600664e2744279a279027ae26a426ba26b61618280411106e497000000e780801c0000197186fca2f8a6f4caf0ceecd2e8d6e4dae0b2891306000232f80d46230cc10203b4090202e002e82af02ef461c003b589026307051083b409009305f5ff8e058d8113891500a10493058003330ab5026104854a17050000130b458a906001caa276027583b584ff946e829665ed08482ad803058401230ca1024c4803b509012eda033684ff0c6001ce631756019205aa95906563046601014621a08c618c61054632e02ee4033684fe833504ff01ce631756019205aa95906563046601014621a08c618c61054632e82eec0c6492052e95106508618a85029649e5c104130a8afc13048403e31b0af6b1a003ba890163080a0483b4090103b409001305faff12051181130915002104a104120a106001caa2760275833584ff946e829639e1906003b584ff8a8502960ded4104411ac104e31e0afc03b589006368a9002da0014903b589006371a90203b5090012092a99a27602758335090003368900946e829619c1054511a00145e6704674a6740679e669466aa66a066b09618280907588711c6e9755ffff938575a12d468287907588711c6e9755ffff938505a139468287411106e497000000e78080010000411106e497000000e780a0000000411106e497b0ffffe780c0170000757106e5014730012948bd4821a89306f6ff13d547009a92a30f56fe0507368663fcf800aa879372f50013030003e3e002ff13037005e1bf13050008198d130610086370c5021755ffff9307a59e09462e85be8597000000e7800082aa60496182809305000897000000e78040660000757106e522e1a6fccaf8cef4d2f0d6ecdae8dee4e2e066fc6af86ef432892e8a014c814c81499715010003bb45d09715010083bb45d09715010083b445d000690c612ef008652aec13058a002ae01755ffff1305c5952ae8294d22e40da03305b6000345f5ff5915133515002300a4006265146d02758296ee8c6311051213f5f90f631b051063758901e9a8636c890d33058941b3058a014146637fc50063022c0d81463386d50003460600630da6098506e319d5fe75a013867500937686ff3386b640ad8e93b6160013371600d98ea1c20146930605ff02676297b387c5009c6313c4f7ffa58fda9733747401e18f8defb307c7009c6313c4f7ffa58fda9733747401e18f95e34106e3f9c6fc31a83387d500034707006307a7038506e319d6fe930605ffe3f9c6fa6304c5062264b386c50083c606006386a6010506e319c5fe05a0b286e296138c1600e3f026f5d29603c50600e31ba5f38149e28de28a39a04a8c8549e68dca8a63872c030345040001c96265146d11460275c265829611ed33869a41b3059a01e39a9aed0145f1bd4a8c2264f9b7014511a00545aa600a64e6744679a679067ae66a466ba66b066ce27c427da27d49618280411106e41b8605009306000802c26376d6002302b100054671a01bd6b50019ee13d665001366060c2302c10093f5f50393850508a302b1000946ada01bd6050115e613d6c5001366060e2302c10013964503699213060608a302c10093f5f503938505082303b1000d462da81396b50275921306060f2302c1001396e502699213060608a302c100139645036992130606082303c10093f5f50393850508a303b10011464c0097000000e780e0d9a26041018280397106fc907594712ae032f836f4886d906994658c612af032ec36e82ee41745ffff9305c57f0a85300097000000e780a0b2e27021618280086117030000670063d5411106e408611b8605009306000802c26376d6002302b100054671a01bd6b50019ee13d665001366060c2302c10093f5f50393850508a302b1000946ada01bd6050115e613d6c5001366060e2302c10013964503699213060608a302c10093f5f503938505082303b1000d462da81396b50275921306060f2302c1001396e502699213060608a302c100139645036992130606082303c10093f5f50393850508a303b10011464c0097000000e78060caa26041018280397106fc90759471986d32f836f43af0906994658c61086132ec36e82ee42ae01745ffff930525700a85300097000000e78000a3e27021618280357106ed22e926e54ae1cefcd2f8d6f42a840345050109c5833a04008544d5a0b2892e89033a840003654a03833a04009375450091e93336500163880a021745ffff9305855d35a063960a0483358a0203350a02946d9745ffff9385255c094682961dc5814a854469a81745ffff9305055b83368a0203350a02946e05068296854441e103b689014a85d28502968da803254a038544a303910283350a0203368a022ee432e8930571022eec83250a0303068a0383360a0003378a0083370a0103388a01aaceaecc2300c10636f43af83efcc2e02800aae403b689011745ffff1305c54faae82c104a85029619e9c6652665946d9745ffff9385055209468296aa8423089400850a233054012285ea604a64aa640a69e679467aa67a0d618280357106ed22e926e54ae1cefcd2f8d6f42a8403458500854a854419cd23049400a30454012285ea604a64aa640a69e679467aa67a0d6182803289ae89033a040003654a03834594001376450005e691cd83358a0203350a02946d9745ffff9385c54909468296854455f94e85d2850299aa846db785e183358a0203350a02946d9745ffff9385c54705468544829659f503254a038544a303910283350a0203368a022ee432e8930571022eec83250a0303068a0383360a0003378a0083370a0103388a01aaceaecc2300c10636f43af83efcc2e02800aae41745ffff1305053eaae82c104e85029915f9c6652665946d9745ffff9385454009468296aa8439bf397106fc22f826f44af02a841c7508719c6f3a89b684829722e8230ca10002e4a30c01002800a6854a8697000000e78060db22658345810139c50544b9e5834591017d1513351500c264b335b0006d8d05c103c54403118901ed8c748870946d9745ffff9385b53905460544829611ed8c748870946d9745ffff93856532054682962a8419a03334b0002285e2704274a274027921618280411106e497000000e78040920000757106e5014730012948bd4831a89306f6ff9377f50f13d547009a92a30f56fe0507368663fbf8001373f50093020003e36f03fd93027003d9bf13050008198d130610086370c5021745ffff9307053109462e85be8597f0ffffe7806014aa60496182809305000897000000e780a0f80000757106e5014730012948bd4831a89306f6ff9377f50f13d547009a92a30f56fe0507368663fbf8001373f50093020003e36f03fd93027005d9bf13050008198d130610086370c5021745ffff9307e52909462e85be8597f0ffffe780400daa60496182809305000897000000e78080f100001745ffff9306e53609462e85b68517f3ffff6700432e397106fc22f826f42e848c752ae40870946d9745ffff9385e5364546829622ec2300a10202e8a30001021745ffff1306653308082c0097000000e780a0c042658345010239c50544b9e5834511027d1513351500e264b335b0006d8d05c103c54403118901ed8c748870946d9745ffff9385f51e05460544829611ed8c748870946d9745ffff9385a517054682962a8419a03334b0002285e2704274a27421618280757106e5014730012948bd4821a89306f6ff13d547009a92a30f56fe0507368663fcf800aa879372f50013030003e3e002ff13037003e1bf13050008198d130610086370c5021745ffff9307651709462e85be8597f0ffffe780c0faaa60496182809305000897000000e78000df0000797106f422f026ec4ae84ee42a8404690865ae893309b640058d6363250308602695ce854a8697f00000e78060dfca9404e8a2700274e2644269a269456182802285a6854a8697000000e780c0000468f9b75d7186e4a2e026fc2e966368b6042a8408659314150063639600b284a14563e39500a14493c5f4fffd9119c5106032f0054632f42af811a002f428001410268697000000e780e003a265426581cdfd55fe158505630ab50009ed97b0ffffe780408a000008e004e4a6600664e27461618280626597b0ffffe78000880000011106ec22e826e44ae03289aa8499cd2e84886605c18c6a91cd88624a8697b0ffffe780808405e180e419a023b40400854521a8630409024a85a28597b0ffffe780a08175d1814588e423b824018ce0e2604264a264026905618280228565f5e1b703e6450308619376060191ea1376060209ee0345050017f3ffff670063d00305050017030000670023d10305050017030000670043c903e6450308619376060189ea1376060219ea086117f3ffff670023cd086117f3ffff67006359086117030000670003e0411106e422e02a8411c96347040289c9228597a0ffffe780407909a8054501a88545228597a0ffffe780a07619c9a285a26002644101828097a0ffffe78000780000228597a0ffffe780a07600005d7186e4a2e026fc4af84ef452f0ae898c750461006903b50902946d9745ffff938525f00546054982964ee42308a100a308010005c417050000930965f1138a140026ec28002c084e8697000000e780e0a17d14d28465f40345010101ed22650c750871946d9745ffff9385f5ef054682962a894a85a6600664e2744279a279027a61618280797106f422f026ec4ae84ee42a8904690865058d2e84636fb50283390900894533859900636cb4007d148145228697f00000e78040aba2943385990023000500850423389900a2700274e2644269a269456182804a85a685228697000000e780e0008334090155bf5d7186e4a2e026fc2e966368b6042a8408659314150063639600b284a14563e39500a14493c5f4fffd9119c5106032f0054632f42af811a002f428001410268697000000e780e003a265426581cdfd55fe158505630ab50009ed97a0ffffe7802062000008e004e4a6600664e27461618280626597a0ffffe780e05f0000011106ec22e826e43284aa8499cd88660dc18c6a99cd8862228697a0ffffe780a05c19ed85458ce431a823b40400854511a88545228597a0ffffe780e0597dd1814588e480e88ce0e2604264a26405618280411106e422e02a8408617d1508e005e90c70086c8c6182950870086511c5086c97a0ffffe780a056087811c5087497a0ffffe780c05508647d1508e409c5a2600264410182802285a2600264410117a3ffff6700c3535d7186e4a2e026fc4af84ef452f056ec83ba0501368a3289aa8963e3da00d28a806108687de1286c7d5610e8637c55010870106c98651c6d4e85b2854a86d286829761a08465306463edc400b386540163ee96082c683307b600636ec7086376d70208700c6c1074147c1c6d0a85268782970345010069e9a26563e8550f286c2ce824e426866367b50eb3b6c400918c33359500558d49e5338554016363950463e7a5080c7c63eca508b3059540639745090c74a6954a85528697f00000e780809623b45901238009000868050508e8a6600664e2744279a279027ae26a616182801745ffff130525e411a81745ffff130585e329a01745ffff1305e5e2f14597f0ffffe780800400001745ffff1305b5d89745ffff9386a5d9c1450a8689a01745ffff1305a5e69305f002d1bf1745ffff1305b5e893052003d9b7528597000000e780e08a00001745ffff1305a5039745ffff938645db9305b0021306710197f0ffffe780801900001745ffff130565dd71b71745ffff130585de9305e00241b7034505000e051746ffff1306c6362a969746ffff9386263b369598751062146188711c6fb6858287411110650c69b29563edc50008611069fd568582637dd60028616369b502410182801745ffff130505aba14535a01745ffff130545cf9745ffff938645d0e145300097f0ffffe780c01000001745ffff130555df9305600297f0ffffe78060f40000797106f422f0aa8502c2280050009146114497000000e78020de0345810011e942656319850203654100a2700274456182801745ffff130545f49745ffff9386e5cb9305b0021306f10197f0ffffe780200a00001745ffff130515dbb54597f0ffffe780e0ed0000411106e497000000e78040f98d4563f7a50009817d15a260410182801745ffff1305e5d8b94597f0ffffe780e0ea0000197186fca2f8a6f4caf0ceecd2e8d6e4dae05efc03bb050003370b00806594692a89130517002330ab0065c95ae409072330eb007dc3b28a36f85af02e8597000000e780a0f29305440063ea850caa892ef4081097000000e780c0f763ffaa02aa84938b1a0013952b002295636e850a2af4081097000000e78040ef2a8a63999b02330544016366850a2ae863f649051745ffff130525ddc1a015452304a900233009005a8597000000e78000c6b1a08a0a33858a002105636285082af4081097000000e78080eab305440163ed8506aa892ee8636e4507338549412aec280097000000e78060e26265c26522662338a9002334b9002330c9005a8597000000e780a0c0e6704674a6740679e669466aa66a066be27b09618280000000001745ffff130545d40da81745ffff1305a5d325a01745ffff130505d339a81745ffff130565d211a81745ffff1305c5d129a01745ffff130525d19305b00297f0ffffe78080d40000797106f422f0906118629465050718e20dcf2a841385460032e4636ad5022ae82e8597000000e78000de2aec280097000000e78020d76265c265226608e80ce410e0a270027445618280000000001745ffff1305e5ca9305b00297f0ffffe78040ce0000397106fc22f826f42a8402e408083000a146a144a28597000000e780c0b70345010105e16265631f9502a264086097000000e780e0b02685e2704274a274216182801745ffff130525cd9745ffff9386c5a49305b0021306710297f0ffffe78000e300001745ffff1305a5b5b94597f0ffffe780c0c60000397106fc22f826f42a84a307010008081306f10085468544a28597000000e78000b0034501010de16265631095048304f100086097000000e78000a92685e2704274a274216182801745ffff130545c59745ffff9386e59c9305b0021306710297f0ffffe78020db00001745ffff130585afb54597f0ffffe780e0be00005d7186e4a2e026fc4af8ae842a898c69054632e002e402e889c90a8597000000e780208f0266426411a001442808a685a28697000000e780a0a6034581011de5027563168504c2652266826688602338b9002334c9002330d900a6600664e27442796161170300006700239e1745ffff130525bb9745ffff9386c5929305b0021306f10297f0ffffe78000d100001745ffff130535a6c94597f0ffffe780c0b40000011106ec22e826e49c692a84637df700b384e74063e3d400b684b306970063ede60263f7d7001545a300a400054531a8998e639dd4028c61ba953285268697e00000e780e03d014504e42300a400e2604264a264056182801745ffff1305658cf14597f0ffffe78000ae00002685b68597f0ffffe780603700005d7186e4a2e026fc4af84ef452f02e8483b905012a896145a14597a0ffffe78020e959c1aa84086888e8086488e4086088e0054a52e402e802ec1314ba002800a28597f0ffffe780007b13050006a14597a0ffffe780c0e531c923304501233445012338050004ed9745ffff938545980cf1a2650cf5c2650cf9e2650cfd23303505233405042338050420ed23340900233839012330a900a6600664e2744279a279027a61618280614519a01305000697a0ffffe780c0e100000c6591c5086117a3ffff670043df8280397106fc22f826f44af09376f60f1307f00f2a89638fe6041b04160002ec02e802e402e0131584036d9113060002098e8a84aa94aa95268597e00000e780002a1375740009c9838504007d563315a6006d8d2380a4008a85130600024a8597e00000e780a027e2704274a274027921618280130600024a858145e2704274a2740279216117e30000670063182a860345050283c605023337d500358d3335a000b306e040558d0de5fd057d06815695c20345060003c70500b337e500398d3335a0003307f040598dfd157d16850665d18280014582805d7186e4a2e026fc4af8ae84806590612a892800a28597e0ffffe78080b30345810019c5426529e109452300a90029a805040dc09305910080e4130610024a8597e00000e780201ca6600664e2744279616182801745ffff1305058cf14597f0ffffe780a08c000097f0ffffe780c0a80000306115ce14610c653337d00093b715007d8f7d1630e115c7106d0c699306050109c683b505227d166dfe0146014723b4060023b00600854614e10ce531a08145b1a8b5ca1869106d83d6a5216374d600ae8621a883b60521a1c603d6852183d7a6210507b685e377f6fe1308160001cf0e083698833708227d1701c783b70722e5bf014811a0b68793050003b305b602b6951ce523380500233c05012e8582801735ffff1305457d9305b00297f0ffffe780a08000001735ffff1305e57bedb7411106e413050022c14597a0ffffe78000bd01c5a260410182801305002297a0ffffe780c0bd0000411106e413050028c14597a0ffffe78080ba01c5a260410182801305002897a0ffffe78040bb00001d7186eca2e8a6e4cae04efc52f856f45af05eec62e866e46ae03e893a8ab689b28aae8b2a84035ca52193841500139b55002a9b139d4500b30cbc40637b9c00130600025a85d68597e00000e780800381a013955400229513965c00da8597e00000e7800047130600025a85d68597e00000e780200113050416b305a50113964400329513964c0097e00000e7806044930a1c00229d23344d1723303d1793092c00130a042213852b00139b3400637c3501b3056a010e05529513963c0097e00000e78000415a9a23302a01231d542163f434038e0ba29b13858b22b305804109461461239c9620850423b88620b38695002105e397c6fee6604664a6640669e279427aa27a027be26b426ca26c026d256182800358a5212e86814593125800aa929303f5011303f601054e63055504938815001305050201579a869e8715cf83ce060003c6070033bfce0033c6ce00b33ec0003306e0413366d601fd17fd16050771de1376f60f631ac60193830302c685e31f55fac28511a0014e72858280457186e7a2e326ff4afb4ef752f356ef5aeb5ee762e3e6feeafaeef62e8a83bb050083b90501b28a2a8b03d9ab21139559005e9583459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18d2ef483451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2ef083459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2eec83451500034605008346250003473500a205d18dc2066207d98ed58d034655008346450003476500834775002206558e4207e2075d8f598e0216d18d2ee8938c190093955c00de9513c6f9ff330426011316540097e00000e780c02093850b16139549002e950465033c050013964c00b2951316440097e00000e780a01e7d3913150903239d2b21033a8a0041919545637bb51a2819de8552869760ffffe780a0736a7556e026e405cd85456317b5068001080113068003a28597e00000e78080d56a65aa750355a52183d5a5212e950505b1456376b50408180c01014605a88001a80013068003a28597e00000e78080d20675c6750355a52183d5a5212e950505b1456372b5040818ac000546ce8697000000e780604899a80e65ae650da0081a13068003a28597e00000e780a0ce081a854597000000e780c0153665d6652af82efccee025a0081a13068003a28597e00000e78020cc081a854597000000e7802072766596752af82efce6e0c27b627a03b60b21866971c613041a00930a010c914c314d954d05498354a62163eb9c0a2819b28522869760ffffe780c0636a751dcd631b2509a81913068003d68597e00000e78020c6526592750355a52183d5a5212e950505636ea503b3859d40a81997000000e780e00b01465df69da0a81913068003d68597e00000e780a0c2526592750355a52183d5a5212e9505056373a503081a13068003d68597e00000e78060c0081a97100000e78080932a862e8425f605a0b3859d40a81997000000e7802065014631fa31a089e4054582652380a500a264227582756266c266233cab002338bb002334cb002330db0023308b0323349b0223387b03233c4b0323303b05be601e64fa745a79ba791a7afa6a5a6bba6b1a6cf67c567db67d79618280317106fd22f926f54af14eed52e956e55ae1defce2f8e6f4eaf0eeec6383052a2e892a8a833b850183d5ab21338425012d45636e85282ef4033b8a020355ab21636e252933052541239d8b202ae4231dab20930af9ff93945a0093090b1613954a002ae84e9583350a01833d0a00106532f008612aec139555006e959205ae9d83459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18daee483451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18daee083459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2efc83451500034605008346250003473500a205d18dc206620703465500d98ecd8e83454500220603476500834775004d8e268cb3059b004207e2075d8f598e0216558e32f81306000297e00000e780e0e403bd0d1683bc8d16626523b0ad16027523b4ad16a28da274139554005e950c181306000297e00000e780409d13840b16139544002295233495018504b3859d402330a501639cba10139554005e95da85628697e00000e780609a139544002295ce85426697e00000e780409993155900da95226c13165c005a8597e00000e780c0dc93154900ce9513164c004e8597e00000e78080db83350a0203350a03adcd79c113040b22139534005e951305052293193900a2854e8697e00000e7800094b305340113163c002106228597e00000e780a0d7a27c63f0bc038e0cde9c13858c220c61239c9520850423b875217d192105e31809fe7d556301ac020145050c0c601306150023b86521239ca52021043285e317ccfe11a039e5ea704a74aa740a79ea694a6aaa6a0a6be67b467ca67c067de66d296182801735ffff13050516ed4505a81735ffff1305151f930520030da01735ffff1305552111a81735ffff1305f50d29a01735ffff1305751a9305800297e0ffffe780c0fa0000317106fd22f926f54af14eed52e956e55ae1defce2f8e6f4eaf0eeec806d035da4216a8701c698750357a721636cd72832f036f42af883ba850203dcaa21930b1d0033868b012d456365c528846188652ae803b9050188712aec03dba42132e4231dc42013155900269583459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18daee883451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18daee483459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18daee083451500034605008346250003473500a205d18dc2066207d98ed58d034655008346450003476500834775002206558e4207e2075d8f598e0216d18d2efc930d190093955d00a6959349f9ffda991396590097e00000e78040b513155d0022952c181306000297d00000e780206f13955b00229513165c00d68597d00000e780e06d93850416131549002e95033a0500833c850013964d00b2951396490097e00000e78080b01305041693154d00aa9523b4950123b0450193850a1613964b00329513164c0097d00000e78020699385042213953d002e950e09ca95c1051396390097e00000e78040ac63f06d032699130589220c6113861d0023b89520239cb5212105b28de317cbfe0395a4217d358545239da420426563f3a50413953b0022951305052293850a2213163c00210697d00000e780806222656372ad02050c0e0d229d13058d22de851061231cb6208505233886207d1c2105e3180cfe02759334150056859790ffffe7804010fd1433f57401a2752e95c27580e1626690e588e9ea704a74aa740a79ea694a6aaa6a0a6be67b467ca67c067de66d296182801735ffff1305f5f49305100939a01735ffff130525fd9305a00297e0ffffe78040cc0000717106f522f126ed4ae94ee552e1d6fcdaf8def4e2f0e6eceae8eee4638605262e8b2a890075835ca421e6952d456363b526033c89018354ac2163e46427338d6441231dac212ee4231db42013155b00229513965c00a28597e00000e780a0989309041613154b004e9513964c00ce8597e00000e7802097930b1d00b38a74411305fbff6396aa2293955b00e295139a5a002285528697d00000e780e04f93040c1693954b00a695920a4e85568697d00000e780604e13154d00269583350901833d0900106532ec08612ae8139555006e959205ae9d83459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18d2efc83451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2ef883459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2ef483451500034605008346250003473500a205d18dc20662070346550083474500d98ecd8e22065d8e034765008347750093155d00e2954207e2075d8f598e0216558e32f01306000297e00000e780a08003bd0d1683b48d16426523b0ad16626523b4ad16330544010c101306000297d00000e7806039d69923b4990023b0a9018335090203350903a1c945c1930404220e0b3385640113963c002106a68597d00000e780407b8e0be29b93850b2226855a8697d00000e780203581452265050590609386150023388620231cb620a104b685e317d5fe11a029e9aa700a74ea644a69aa690a6ae67a467ba67b067ce66c466da66d4d6182801735ffff1305c5baed4515a81735ffff1305b5bb930530031da01735ffff130505be9305700221a81735ffff130575b229a01735ffff1305f5be9305800297e0ffffe780409f0000357106ed22e926e54ae1cefcd2f8d6f4daf0deece2e8e6e4eae06efc033a850183398502835aaa2103dba92113841a0033066401ad4563e1c526033d0500833c050108652ae8035cad2132e4231dca2013955c006a9583459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18d2ef883451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2ef483459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2ef083451500034605008346250003473500a205d18dc2066207d98ed58d034655008346450003476500834775002206558e4207e2075d8f598e0216d18d2eec93841c0093955400ea9593cdfcffe29d13965d0097d00000e780005b13955a0052952c081306000297d00000e780e01413155400529513165b00ce8597d00000e780a01393050d1613954c002e9503390500833b850013964400b29513964d0097d00000e780405613050a1693954a00aa9523b4750123b025019385091613164400329513164b0097d00000e780e00e93050d22139534002e958e0ce695c10513963d0097d00000e780005263f08403ea9c13858c220c611386140023b8a521239c95202105b284e317ccfe0315ad217d358545231dad20c26463f29504131534005295130505229385092213163b00210697d00000e7804008226563f1aa02050b8e0ad29a13858a220c61239c8520050423b845217d1b2105e3180bfe4e859790ffffe78080b66a85a685ea604a64aa640a69e679467aa67a067be66b466ca66c066de27d0d6182801735ffff130545a59305a00297d0ffffe78060740000411106e413058072a1459790ffffe78060b101c5a26041018280130580729790ffffe78020b20000411106e413058078a1459790ffffe780e0ae01c5a26041018280130580789790ffffe780a0af00001d7186eca2e8a6e4cae04efc52f856f45af05eec62e866e43a89b689328a2e8b2a84835b655b1305855b938415009605da95b30ab500338c6b4163fb9b00130610025685d28597d00000e78000f8a9a09395540026952e9513165c006296d68597d00000e780403b130610025685d28597d00000e78060f51305840013064008b305cb02aa95b386c40236953306cc0297d00000e7804038138a1b00130540083305ab022295210513064008ce8597d00000e78080f193892b00930a847213052b00939c3400637c3501b3859a010e05569513163c0097d00000e780e033e69a23b02a01231b445b63f334030e0b229b13050b73b305704109461461239a965a850480e2b38695002105e398c6fee6604664a6640669e279427aa27a027be26b426ca26c25618280397106fc22f826f44af04eec52e856e48359655b2e8a9305855b93945900ce947d54054995c4938a1502528597f0ffffe78060c29384f4fd1375f50f0504d685e30225ff9305f00f6305b500014911a04e844a85a285e2704274a2740279e269426aa26a21618280130101ce233c1130233881302334913023302131233c312f2338412f2334512f2330612f233c712d2338812d2334912d2330a12d233cb12b2e8c83bb050003bb05013289aa8903da6b5b13848b5b13155b005a95b30ca400a80b13061002e68597d00000e78060dd930a1b0093955a005694a2951345fbffb3044501139654002696668597d00000e7800020930c400833059b033384ab00130d84001305911f13064008ea8597d00000e78000d99305c408338694036a8597d00000e780c01c1b05faff239bab5a033a8c004215135405032811ac0b1306500a97d00000e780c0d50a852c111306500a97d00000e780c0d41545637da41a2811de85528697000000e78060202a7505cd85456317b5060019081313068003a28597d00000e780c0d17a75be650355655b83d5655b2e950505b1456376b504880a0c13014605a80019a81213068003a28597d00000e780c0ce1a65da650355655b83d5655b2e950505b1456372b504880aac120546da8697000000e780004ca9a84a75ea750da0a80b13068003a28597d00000e780e0caa80b854597000000e780601d5e75fe75aaeaaeeedaf235a0a80b13068003a28597d00000e78060c8a80b854597000000e780a06b0335012083358120aaeaaeeed6f2d66b766a03b60b00167b69ca93041a00930a010b914d314c954c054d0354665b63ee8d0a2811b285268697000000e78080102a7529c1631fa509080513068003d68597d00000e78020c2033581298335812a0355655b83d5655b2e95050563608505b3858c40080597000000e780001301464df6a5a0080513068003d68597d00000e78060be033581298335812a0355655b83d5655b2e95050563738503a80b13068003d68597d00000e780e0bba80b97100000e78020882a86ae8425f239a8b3858c40080597000000e780e05d014631f629a001e405452300a9008a851306500a4e8597d00000e78000b823b4790b23b8490b23bc690b833081310334013183348130033901308339812f033a012f833a812e033b012e833b812d033c012d833c812c033d012c833d812b13010132828094619dc683d7455b130816009dc71387f7ff93173700b69783b787722330050014e52338050118ed1cf110f50cf92da00ce510e989450ce1828003d7665b19cf03b7067385471ce114e523380501233c05000cf110f518f910fd828097d0ffffe780803c0000130101d92334112623308126233c9124233821252334312523304125233c5123233861232334712323308123233c91212338a1212334b121638505242e89aa8b033d850103546d5bb304b4002d456360952422ec83bc8b0203d56c5b63602525330a2541231b9d5a239b4c5b930df9ff93898c5b13955d006e952ae4338ba900938a8c0013044008b3858d022ee8d69528101306400897d00000e78060a303b50b0183b50b0013165500b386a500369626f09304865b330585022e95130c8500081913061002a68597d00000e78040a0130610022685da8597d00000e78020e49304110d130640082685e28597d00000e780009e2c1013064008628597d00000e780009da80a0c191306100297d00000e780009c080313064008a68597d00000e780009b130b8d5b626c13155c00b3058b012e95ac0a1306100297d00000e780209993048d0033058c0226950c031306400897d00000e780a09713041c000275018d6392ad1413155400229b5a95ce85226697d00000e780a095130b4008330564032695d685426697d00000e7804094131559004a95b385a90013165a0052964e8597d00000e78080d7b3056903d69533066a03568597d00000e78040d683b50b0203b50b03c1c165c5d28a93848c72131534006a951305857293193900a6854e8697d00000e780a08eb385340113163a002106268597d00000e78040d202756371ac02131a3c006a9a13050a730c61239a855a050423b0a5017d192105e31809fe7d556382aa02814513851a0090609386150023309601231ab65aa104b685e317d5fe11a02de58330812603340126833481250339012583398124033a0124833a8123033b0123833b8122033c0122833c8121033d0121833d81201301012782801725ffff1305a50eed4505a81725ffff1305b517930520030da01725ffff1305f51911a81725ffff1305950629a01725ffff130515139305800297d0ffffe78060f30000697106f622f226ee4aea4ee652e2d6fddaf9def5e2f1e6edeae9eee583bd850103dc6d5b628701c698750357675b636ad71e32f036f42af883ba850283dc6a5b130b1c0033069b012d456363c51e846188652ae888712aec83b9050183db645b32e4239bcd5a1384845b139559004e95330da400880013061002ea8597c00000e780a07813891900931559004a94a29513caf9ff5e9a52fc13165a0052966a8597d00000e78040bb13848d5b13155c00b30584012e958c001306100297c00000e780a07493858a5b13155b005a94229513965c00669697c00000e7800073130d40083385a9033384a400628a5a8c668bd68c930a8400880013064008d68597c00000e78080709305c40862753306a5035685e68ada8c628b97d00000e780c0b313848d003305aa0322958c001306400897c00000e780606d93858a003305ac0322953386ac0397c00000e780006c93858472131539002e958e09ce95c10562760e0697d00000e78020af637f7901a699138509730c611306190084e1239a255b21053289e398cbfe0395645b7d358545239ba45a426563f4a50413153b006e951305857293858a7213963c00210697c00000e780806522656373aa02850c131c3a006e9c13050c73da851061231ab65a85052330b601fd1c2105e3980cfe02751334150056859780ffffe78020137d1433756401a2752e95c27523b0b501626690e588e9b2701274f2645269b269126aee7a4e7bae7b0e7cee6c4e6dae6d556182801725ffff1305b5f79305100939a01725ffff1305e5ff9305a00297d0ffffe78000cf0000130101d92334112623308126233c9124233821252334312523304125233c5123233861232334712323308123233c91212338a1212334b121638705202e8caa8b0075035d645bea952d456364b52003bb8b01835a6b5b63e58a21338a8a41231b4b5b2ee8231bb45a1309845b13155c0062954a9513165d006a96ca8597d00000e780209993098400930c400833059c034e9533069d03ce8597d00000e7806097930d1a00b384ba411305fcff6391a41cda8a130b8b5b93955d003305bb01aa95139554003306950032f04a8597c00000e780404f56e4a10ab3859d03d6953386940332ec4e8597c00000e780a04d13155a00529b2a9bb3059a03d69528101306400897c00000e780e04b03b50b0183b50b0013165500b386a50036969304865b330595032e95930c8500081913061002a68597c00000e780e048130610022685da8597d00000e780c08c9304110d130640082685e68597c00000e780a0462c1013064008668597c00000e780a045a80a0c191306100297c00000e780a044080313064008a68597c00000e780a04302754a95ac0a1306100297c00000e780804262654e950c031306400897c00000e780604183b50b0203b50b03a1c955cd930484720e0c3385840113163d002106a68597d00000e780e0838e0d2265aa9d93858d722685628697c00000e780a03d81454265050590609386150000e2231ab65aa104b685e318d5fe11a03de58330812603340126833481250339012583398124033a0124833a8123033b0123833b8122033c0122833c8121033d0121833d81201301012782801725ffff1305a5c1ed4515a81725ffff130595c2930530031da01725ffff1305e5c49305700221a81725ffff130555b929a01725ffff1305d5c59305800297d0ffffe78020a600006d7106e622e2a6fdcaf9cef5d2f1d6eddae9dee5e2e166fd6af96ef5033a850183398502035b6a5b83db695b13041b0033067401ad4563ebc51a833c05000c652eec833d050103dd6c5b32e0231bca5a13898c5b13955d006e95b30aa900081013061002d68597c00000e780c02c93841d00939554002699ca9513c9fdff6a99131659004a96568597c00000e780806f930a8a5b13155b00b3856a012e950c101306100297c00000e780e0289385895b13155400a29a569513965b005e9697c00000e7804027130c400833858d03b38aac005ee4ce8b93898a00081013064008ce8597c00000e78000259385ca08330689034e8597c00000e780c06893098a005ae833058b034e950c101306400897c00000e7804022de8a93858b00a26b330584034e9533868b0397c00000e780a02093858c72139534002e958e0dee95c1051316390097c00000e780c06363f0a403e69d13850d730c611386140023b09501239a955a2105b284e317cdfe03956c5b7d358545239bac5ae264426b63f295041315340052951305857293858a7213963b00210697c00000e780e01902656371ab02850b0e0b529b13050b730c61239a855a050423b04501fd1b2105e3980bfe56859780ffffe78020c86685a685b2601264ee744e79ae790e7aee6a4e6bae6b0e6cea7c4a7daa7d516182801725ffff1305e5b69305a00297d0ffffe78000860000130101dc233c1122233881222334912223302123233c3121233841212334512123306121deffe2fbe6f7eaf3eeefd54bae8a63f575052a8c094563e9aa0005466285d68597300000e78060e98330812303340123833481220339012283398121033a0121833a8120033b0120fe7b5e7cbe7c1e7dfe6d130101248280b68cb2892afc930d7113054d0545aae856f8627c1b850c0019e16f20f00613751d0019e16f10b07d466813db2a0013171b00b308670113051003637955231303fbff93021b0013166b00629603459601834586018346a6018347b60122054d8dc206e207dd8e558d8345d6018346c6018347e6018344f601a205d58dc207e204c58fdd8d82154d8d2af90345160183450601834626018347360122054d8dc206e207dd8e558d83455601834646018347660183447601a205d58dc207e204c58fdd8d82154d8d2af503459600834586008346a6008347b60022054d8dc206e2078345d6008344c600dd8e558da205cd8c8346e6008347f60093156300e295c206e207dd8ec58e8216558d2af1034516008346060083472600834436002205558dc207e204c58f5d8d83465600834746008344660003467600a206dd8ec2046206458e558e0216518d2aed03c5950103c6850183c6a50183c7b5012205518dc206e207dd8e558d03c6d50183c6c50183c7e50183c4f5012206558ec207e204c58f5d8e0216518d2afa03c5150103c6050183c6250183c735012205518dc206e207dd8e558d03c6550183c6450183c7650183c475012206558ec207e204c58f5d8e0216518d2af603c5950003c6850083c6a50083c7b5002205518dc206e207dd8e558d03c6d50083c6c50083c7e50083c4f5002206558ec207e204c58f5d8e0216518d2af203c5150003c6050083c6250083c735002205518dc206e207dd8e558d03c6550083c6450083c7650083c575002206558ec207e205dd8dd18d82154d8d2aee01559305710b6e8605c583c60500834706007d16fd150505e388f6feb3b3f60063f9f6009a875a8331a081436f10c0168143da8713956200629503469501834685018344a5010344b5012206558ec2046204458c418e8346d5018344c5010344e5018345f501a206c58e4204e205c18dd58d8215d18d2ef983451501034605018346250183443501a205d18dc206e204c58ed58d034655018346450183446501034475012206558ec2046204458c418e0216d18d2ef583459500034685008346a5008344b500a205d18dc206e2040346d5000344c500c58ed58d2206518c8346e5008344f500139667006296c206e204c58ec18e8216d58d2ef183451500834605008344250003443500a205d58dc2046204458cc18d83465500834445000344650003457500a206c58e42046205418d558d02154d8d2aed03459601834586018346a6018344b60122054d8dc206e204c58e558d8345d6018346c6018344e6010344f601a205d58dc2046204458cc18d82154d8d2afa0345160183450601834626018344360122054d8dc206e204c58e558d83455601834646018344660103447601a205d58dc2046204458cc18d82154d8d2af603459600834586008346a6008344b60022054d8dc206e204c58e558d8345d6008346c6008344e6000344f600a205d58dc2046204458cc18d82154d8d2af20345160083450600834626008344360022054d8dc206e204c58e558d83455600834646008344660003467600a205d58dc2046206458ed18d82154d8d2aee01551306710b130471130dc183440600834604007d147d160505e388d4fe63e3d400be8233b5d400aa93968713956700629583459501034685018346a5018344b501a205d18dc206e204c58ed58d0346d5018346c5018344e5010344f5012206558ec2046204458c418e0216d18d2ef983451501034605018346250183443501a205d18dc206e204c58ed58d034655018346450183446501034475012206558ec2046204458c418e0216d18d2ef583459500034685008346a5008344b500a205d18dc206e2040346d5000344c500c58ed58d2206518c8346e5008344f500131663006296c206e204c58ec18e8216d58d2ef183451500834605008344250003443500a205d58dc2046204458cc18d83465500834445000344650003457500a206c58e42046205418d558d02154d8d2aed03459601834586018346a6018344b60122054d8dc206e204c58e558d8345d6018346c6018344e6010344f601a205d58dc2046204458cc18d82154d8d2afa0345160183450601834626018344360122054d8dc206e204c58e558d83455601834646018344660103447601a205d58dc2046204458cc18d82154d8d2af603459600834586008346a6008344b60022054d8dc206e204c58e558d8345d6008346c6008344e6000344f600a205d58dc2046204458cc18d82154d8d2af20345160083450600834626008344360022054d8dc206e204c58e558d83455600834646008344660003467600a205d58dc2046206458ed18d82154d8d2aee01551306710b9304711315c10344060083c60400fd147d160505e308d4fe6363d4003e833335d400aa931a8b11a03e8b9304f7ff9362170013156700629583459501034685018346a5018347b501a205d18dc206e207dd8ed58d0346d5018346c5018347e5010344f5012206558ec2076204c18f5d8e0216d18d2ef983451501034605018346250183473501a205d18dc206e207dd8ed58d034655018346450183476501034475012206558ec2076204c18f5d8e0216d18d2ef583459500034685008346a5008347b500a205d18dc206e2070346d5000344c500dd8ed58d2206518c8346e5008347f500139664006296c206e207dd8ec18e8216d58d2ef183451500834605008347250003443500a205d58dc2076204c18fdd8d83465500834745000344650003457500a206dd8e42046205418d558d02154d8d2aed03459601834586018346a6018347b60122054d8dc206e207dd8e558d8345d6018346c6018347e6010344f601a205d58dc2076204c18fdd8d82154d8d2afa0345160183450601834626018347360122054d8dc206e207dd8e558d83455601834646018347660103447601a205d58dc2076204c18fdd8d82154d8d2af603459600834586008346a6008347b60022054d8dc206e207dd8e558d8345d6008346c6008347e6000344f600a205d58dc2076204c18fdd8d82154d8d2af20345160083450600834626008347360022054d8dc206e207dd8e558d83455600834646008347660003467600a205d58dc20762065d8ed18d82154d8d2aee01551306710b9306711315c18347060003c40600fd167d160505e38887fe33b58700aa9363f58700a686ba8411a0ba8613956200629583459501034685010347a5018347b501a205d18d4207e2075d8fd98d0346d5010347c5018347e5010344f5012206598ec2076204c18f5d8e0216d18d2ef983451501034605010347250183473501a205d18d4207e2075d8fd98d034655010347450183476501034475012206598ec2076204c18f5d8e0216d18d2ef583459500034685000347a5008347b500a205d18d4207e2070346d5000344c5005d8fd98d2206518c0347e5008347f5001396660062964207e2075d8f418f0217d98d2ef183451500034705008347250003443500a205d98dc2076204c18fdd8d0347550083474500034465000345750022075d8f42046205418d598d02154d8d2aed03459601834586010347a6018347b60122054d8d4207e2075d8f598d8345d6010347c6018347e6010344f601a205d98dc2076204c18fdd8d82154d8d2afa0345160183450601034726018347360122054d8d4207e2075d8f598d83455601034746018347660103447601a205d98dc2076204c18fdd8d82154d8d2af603459600834586000347a6008347b60022054d8d4207e2075d8f598d8345d6000347c6008347e6000344f600a205d98dc2076204c18fdd8d82154d8d2af20345160083450600034726008347360022054d8d4207e2075d8f598d83455600034746008347660003467600a205d98dc20762065d8ed18d82154d8d2aee01551306710b130771130dc103440600834707007d177d160505e308f4fe6363f400b6823335f400aa93968613956600629583459501034685010347a5018347b501a205d18d4207e2075d8fd98d0346d5010347c5018347e5010344f5012206598ec2076204c18f5d8e0216d18d2ef983451501034605010347250183473501a205d18d4207e2075d8fd98d034655010347450183476501034475012206598ec2076204c18f5d8e0216d18d2ef583459500034685000347a5008347b500a205d18d4207e2070346d5000344c5005d8fd98d2206518c0347e5008347f5001396640062964207e2075d8f418f0217d98d2ef183451500034705008347250003443500a205d98dc2076204c18fdd8d0347550083474500034465000345750022075d8f42046205418d598d02154d8d2aed03459601834586010347a6018347b60122054d8d4207e2075d8f598d8345d6010347c6018347e6010344f601a205d98dc2076204c18fdd8d82154d8d2afa0345160183450601034726018347360122054d8d4207e2075d8f598d83455601034746018347660103447601a205d98dc2076204c18fdd8d82154d8d2af603459600834586000347a6008347b60022054d8d4207e2075d8f598d8345d6000347c6008347e6000344f600a205d98dc2076204c18fdd8d82154d8d2af20345160083450600034726008347360022054d8d4207e2075d8f598d83455600034746008347660003467600a205d98dc20762065d8ed18d82154d8d2aee01551306710b1307711315c183470600034407007d177d160505e38887fe63e38700b68433b58700aa93268711a036871383f8ff9382180013956800629583459501034685018346a5018347b501a205d18dc206e207dd8ed58d0346d5018346c5018347e5018344f5012206558ec207e204c58f5d8e0216d18d2ef983451501034605018346250183473501a205d18dc206e207dd8ed58d034655018346450183476501834475012206558ec207e204c58f5d8e0216d18d2ef583459500034685008346a5008347b500a205d18dc206e2070346d5008344c500dd8ed58d2206d18c8346e5008347f500131663006296c206e207dd8ec58e8216d58d2ef183451500834605008347250083443500a205d58dc207e204c58fdd8d83465500834745008344650003457500a206dd8ec2046205458d558d02154d8d2aed03459601834586018346a6018347b60122054d8dc206e207dd8e558d8345d6018346c6018347e6018344f601a205d58dc207e204c58fdd8d82154d8d2afa0345160183450601834626018347360122054d8dc206e207dd8e558d83455601834646018347660183447601a205d58dc207e204c58fdd8d82154d8d2af603459600834586008346a6008347b60022054d8dc206e207dd8e558d8345d6008346c6008347e6008344f600a205d58dc207e204c58fdd8d82154d8d2af20345160083450600834626008347360022054d8dc206e207dd8e558d83455600834646008347660003467600a205d58dc20762065d8ed18d82154d8d2aee01551306710b9304711315c18346060083c70400fd147d160505e388f6fe33b5f600aa9363f5f6001a86468311a0468613956200629583459501834685018347a5018344b501a205d58dc207e204c58fdd8d8346d5018347c5018344e5010344f501a206dd8ec2046204458cc18e8216d58d2ef983451501834605018347250183443501a205d58dc207e204c58fdd8d83465501834745018344650103447501a206dd8ec2046204458cc18e8216d58d2ef583459500834685008347a5008344b500a205d58dc207e2048346d5000344c500c58fdd8da206c18e8347e5000344f50093146600e294c2076204c18fdd8e8216d58d2ef183451500834605008347250003443500a205d58dc2076204c18fdd8d83465500834745000344650003457500a206dd8e42046205418d558d02154d8d2aed03c5940183c5840183c6a40183c7b40122054d8dc206e207dd8e558d83c5d40183c6c40183c7e40103c4f401a205d58dc2076204c18fdd8d82154d8d2afa03c5140183c5040183c6240183c7340122054d8dc206e207dd8e558d83c5540183c6440183c7640103c47401a205d58dc2076204c18fdd8d82154d8d2af603c5940083c5840083c6a40083c7b40022054d8dc206e207dd8e558d83c5d40083c6c40083c7e40003c4f400a205d58dc2076204c18fdd8d82154d8d2af203c5140083c5040083c6240083c7340022054d8dc206e207dd8e558d83c5540083c6440083c7640083c47400a205d58dc207e204c58fdd8d82154d8d2aee01559304710b130471130dc183c70400834604007d14fd140505e388d7fe63e3d700b28233b5d700aa93168613156600629583459501834685018347a5018344b501a205d58dc207e204c58fdd8d8346d5018347c5018344e5010344f501a206dd8ec2046204458cc18e8216d58d2ef983451501834605018347250183443501a205d58dc207e204c58fdd8d83465501834745018344650103447501a206dd8ec2046204458cc18e8216d58d2ef583459500834685008347a5008344b500a205d58dc207e2048346d5000344c500c58fdd8da206c18e8344e5000344f50093176300e297c2046204458cc18e8216d58d2ef183451500834605008344250003443500a205d58dc2046204458cc18d83465500834445000344650003457500a206c58e42046205418d558d02154d8d2aed03c5970183c5870183c6a70183c4b70122054d8dc206e204c58e558d83c5d70183c6c70183c4e70103c4f701a205d58dc2046204458cc18d82154d8d2afa03c5170183c5070183c6270183c4370122054d8dc206e204c58e558d83c5570183c6470183c4670103c47701a205d58dc2046204458cc18d82154d8d2af603c5970083c5870083c6a70083c4b70022054d8dc206e204c58e558d83c5d70083c6c70083c4e70003c4f700a205d58dc2046204458cc18d82154d8d2af203c5170083c5070083c6270083c4370022054d8dc206e204c58e558d83c5570083c6470083c4670083c77700a205d58dc204e207c58fdd8d82154d8d2aee01559307710b9304711315c103c4070083c60400fd14fd170505e308d4fe6363d40032833335d400aa939a8811a0b28813156700629503469501834685018347a5018344b5012206558ec207e204c58f5d8e8346d5018347c5018344e5010344f501a206dd8ec2046204458cc18e8216558e32f9034615018346050183472501834435012206558ec207e204c58f5d8e83465501834745018344650103447501a206dd8ec2046204458cc18e8216558e32f503469500834685008347a5008344b5002206558ec207e2048346d5000344c500c58fd18fa206c18e8344e5000344f50013166b006296c2046204458cc18e8216dd8e36f183461500834705008344250003443500a206dd8ec2046204458cc18e83475500834445000344650003457500a207c58f42046205418d5d8d0215558d2aed03459601834686018347a6018344b6012205558dc207e204c58f5d8d8346d6018347c6018344e6010344f601a206dd8ec2046204458cc18e8216558d2afa034516018346060183472601834436012205558dc207e204c58f5d8d83465601834746018344660103447601a206dd8ec2046204458cc18e8216558d2af603459600834686008347a6008344b6002205558dc207e204c58f5d8d8346d6008347c6008344e6000344f600a206dd8ec2046204458cc18e8216558d2af2034516008346060083472600834436002205558dc207e204c58f5d8d83465600834746008344660003467600a206dd8ec2046206458e558e0216518d2aee01551306710b9306711315c18347060083c40600fd167d160505e38897fe33b59700aa9363f597005a863a8b11a03a8613956800629583469501034785018347a5018344b501a206d98ec207e204c58fdd8e0347d5018347c5018344e5010344f50122075d8fc2046204458c418f0217d98e36f983461501034705018347250183443501a206d98ec207e204c58fdd8e0347550183474501834465010344750122075d8fc2046204458c418f0217d98e36f583469500034785008347a5008344b500a206d98ec207e2040347d5000344c500c58fd58f2207418f8344e5000344f50093166600e296c2046204458c418f02175d8f3af10347150083470500834425000344350022075d8fc2046204458c418f83475500834445000344650003457500a207c58f42046205418d5d8d0215598d2aed03c5960103c7860183c7a60183c4b6012205598dc207e204c58f5d8d03c7d60183c7c60183c4e60103c4f60122075d8fc2046204458c418f0217598d2afa03c5160103c7060183c7260183c436012205598dc207e204c58f5d8d03c7560183c7460183c4660103c4760122075d8fc2046204458c418f0217598d2af603c5960003c7860083c7a60083c4b6002205598dc207e204c58f5d8d03c7d60083c7c60083c4e60003c4f60022075d8fc2046204458c418f0217598d2af203c5160003c7060083c7260083c436002205598dc207e204c58f5d8d03c7560083c7460083c4660083c6760022075d8fc204e206c58ed98e8216558d2aee01559306710b130771130dc183c70600834407007d17fd160505e38897fe63e39700b28833b59700aa93468613156600629583469501034785018347a5018344b501a206d98ec207e204c58fdd8e0347d5018347c5018344e5010344f50122075d8fc2046204458c418f0217d98e36f983461501034705018347250183443501a206d98ec207e204c58fdd8e0347550183474501834465010344750122075d8fc2046204458c418f0217d98e36f583469500034785008347a5008344b500a206d98ec207e2040347d5000344c500c58fd58f2207418f8344e5000344f50093166b00e296c2046204458c418f02175d8f3af10347150083470500834425000344350022075d8fc2046204458c418f83475500834445000344650003457500a207c58f42046205418d5d8d0215598d2aed03c5960103c7860183c7a60183c4b6012205598dc207e204c58f5d8d03c7d60183c7c60183c4e60103c4f60122075d8fc2046204458c418f0217598d2afa03c5160103c7060183c7260183c436012205598dc207e204c58f5d8d03c7560183c7460183c4660103c4760122075d8fc2046204458c418f0217598d2af603c5960003c7860083c7a60083c4b6002205598dc207e204c58f5d8d03c7d60083c7c60083c4e60003c4f60022075d8fc2046204458c418f0217598d2af203c5160003c7060083c7260083c436002205598dc207e204c58f5d8d03c7560083c7460083c4660083c6760022075d8fc204e206c58ed98e8216558d2aee01559306710b130771130dc183c70600834407007d17fd160505e38897fe63f797002d4563f4a356850311a0328b13b513003375a8006319055a13146b00638f095ae3765b63b3048c0003c5990183c5890103c6a90183c6b90122054d8d4206e206558e518d83c5d90103c6c90183c6e90103c7f901a205d18dc2066207d98ed58d82154d8d2af903c5190183c5090103c6290183c6390122054d8d4206e206558e518d83c5590103c6490183c6690103c77901a205d18dc2066207d98ed58d82154d8d2af503c5990083c5890003c6a90083c6b90022054d8d4206e206558e518d83c5d90003c6c90083c6e90003c7f900a205d18dc2066207d98ed58d82154d8d2af103c5190083c5090003c6290083c6390022054d8d4206e206558e518d83c5590003c6490083c6690003c77900a205d18dc2066207d98ed58d82154d8d2aed03c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8d2afa03c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8d2af603c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8d2af203c5140083c5040003c6240083c6340022054d8d4206e206558e518d83c5540003c6440083c6640003c77400a205d18dc2066207d98ed58d82154d8d2aee01559305710b1306711301cd83c60500034706007d16fd150505e388e6fe63e5e63a4e89280a13060004e28597a00000e7804042130600046285a68597b00000e78020862c0a13060004268597a00000e780404093090c04280913060004e28597a00000e780003f0144568b1305fbff6370a414130871139308711b93156400ce954a76aa760a77ea6732fb36f73af33eef03c6950183c6850103c7a50183c7b5012206558e4207e2075d8f598e83c6d50103c7c50183c7e50183c4f501a206d98ec207e204c58fdd8e8216558e32fa03c6150183c6050103c7250183c735012206558e4207e2075d8f598e83c6550103c7450183c7650183c47501a206d98ec207e204c58fdd8e8216558e32f603c6950083c6850003c7a50083c7b5002206558e4207e2075d8f598e83c6d50003c7c50083c7e50083c4f500a206d98ec207e204c58fdd8e8216558e32f203c6150083c6050003c7250083c735002206558e4207e2075d8f598e83c6550003c7450083c7650083c57500a206d98ec207e205dd8dd58d8215d18d2eee81554686c28681cd0347060083c70600fd167d168505e308f7fe6366f7000504e319a4ec2a84637aa4162a8b93146500e2944a75aa750a76ea662afb2ef732f336ef03c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8d2afa03c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8d2af603c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8d2af203c5140083c5040003c6240083c6340022054d8d4206e20683c55400558e498e03c54400a20583c6640003c77400c98d1305fbffc2066207d98ed58d8215d18d2eee81551306711b9306711381cd0347060083c70600fd167d168505e308f7fee365f7ec131a64004e9a280a13060004d28597a00000e7808015130600045285a68597a00000e78060592c0a13060004268597a00000e78080130504a9b3930414002c0913060004628597a00000e7800012e3eb9a10b38a9a409a04269cca8963e47a016fe06f866fe0af80014593d81a0013966a00b304cc00e286130700fcb6873386e4000304060083850700238087002300b6000507850765f70505938404fc93860604e31b15fd134bfbff569b054585b46285d68597200000e780a0c40148fd3c6fe0cf816285d68597200000e78060d8e30305a46fd0fffa627c427a11a0568a13097113130d710be3784b076294280a13060004e28597a00000e7800007130600046285a28597a00000e780e04a2c0a13060004228597a00000e7800005930b0c04930afaffa80813060004e28597a00000e78080030144131564005e9583459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18d2ef983451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2ef583459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2ef183451500034605008346250003473500a205d18dc2066207d98ed58d034655008346450003476500034575002206558e42076205598d518d02154d8d2aed4675a6750676e6662afa2ef632f236ee01559305710b1306711305c183c60500034706007d16fd150505e388e6fe63f6e6000504e31754ed5684d685ae84637bb41213956400629583459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18d2ef983451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2ef583459500034685008346a5000347b500a205d18dc20662070346d500d98ecd8e8345c50022060347e5008347f5004d8e9385f4ff4207e2075d8f598e0216558e32f1034615008346050003472500834735002206558e4207e2075d8f598e83465500034745008347650003457500a206d98ec20762055d8d558d0215518d2aed46752676867666672afa32f636f23aee01556a86ca86e30105ee0347060083c70600fd167d160505e307f7fee376f7ec63ef845a62fc4ef066e852f863e79a5a814a8149014b814d26e43385844022f493156400de951a05338ca50093030008130300082eecae8b130871079302101033057c41135e650063775e0233b56d01b3b55901c98d3305b040137505f872952a8663e46d011e862a83b28389e513531500b303654063856d01639e5929a1aa630503148145130b81095e859308711b03469501834685010347a5018347b5012206558e4207e2075d8f598e8346d5010347c5018347e5010344f501a206d98ec2076204c18fdd8e8216558e32fb034615018346050103472501834735012206558e4207e2075d8f598e83465501034745018347650103447501a206d98ec2076204c18fdd8e8216558e32f703469500834685000347a5008347b5002206558e4207e2075d8f598e8346d5000347c5008347e5000344f500a206d98ec2076204c18fdd8e8216558e32f3034615008346050003472500834735002206558e4207e20783465500034445005d8f598ea206c18e03476500834775002300bb0085054207e2075d8fd98e8216558e32ef0156c686428715c283c7060003440700b3b48700a18f3334f000b3079040c18f7d17fd160506e5d311a0814713b6f7ff329b13050504e39665ec19a0130b8109930d810963925915638c03120145930a8111e2859308711b2380aa00050503c695fd83c685fd03c7a5fd83c7b5fd2206558e4207e2075d8f598e83c6d5fd03c7c5fd83c7e5fd83c4f5fda206d98ec207e204c58fdd8e8216558e32fb03c615fd83c605fd03c725fd83c735fd2206558e4207e2075d8f598e83c655fd03c745fd83c765fd83c475fda206d98ec207e204c58fdd8e8216558e32f703c695fc83c685fc03c7a5fc83c7b5fc2206558e4207e2075d8f598e83c6d5fc03c7c5fc83c7e5fc83c4f5fca206d98ec207e204c58fdd8e8216558e32f303c615fc83c605fc03c725fc83c735fc2206558e4207e2075d8f598e83c645fc03c755fc83c765fc83c475fc938505fc2207d98ec207e204c58fdd8e8216558e32ef0156c686428701ce83c70600034407007d17fd160506e38887fe33b68700b29ae31f75ec19a0930a8111930981113309bb4133853a416363a9002a896309090cf2e09ee49ae803c50d001a05b385ab00280b1306000497a00000e780e0a703ca090003c50d00934cfaff93956c00e2951a05de845e951306000497a00000e780a0a505456315a900ce8b6e8d99a87d1903c51d00138d1d001a053384a4001345faff136505f01a05629513060004a28597a00000e78040a203ca1900938b1900934cfaff93956c00e29513060004228597a00000e78040a07d19ea8dde89e31909fa13956c0062952c0b1306000497a00000e780609e930d1d0093891b001308710793021010a68b4663a663066e33c56d013335a0007d15337565001a05aa9b33c559013335a000b30570407d156d8d1a052a9ce3725ec263f86d0562840345fbff1309fbff1a05b384ab00130404fc280b13060004a68597a00000e780c097130600042685a28597a00000e780a0db2c0b13060004228597a00000e780c0954a8be3ee2dfb91a85e8463f8590503c5faff1389faff1345f5ff1a05b304ac00280b13060004a28597a00000e780c092130600042285a68597a00000e780a0d62c0b13060004268597a00000e780c09013040404ca8ae3ec29fb62653305a4401981a27aaa9aac08130600046274228597a00000e780408ec27463f99a0c139c6a00229c280a13060004a28597a00000e780808c130600042285e28597a00000e78060d02c0a13060004628597a00000e780808a33845441568963e38a0022897d1493090c04d54bc26c930d711363fe8a006275d6850276e68697d0ffffe780a07462f0a28a4e8c11a84e85a2856286e68697d0ffffe7802073627c2275a2653335b50013451500aae813d534003335a900134d150056f862fc827963e47a016fd02ff96fd08ff36285d68597100000e780809d6fd0cff35a85d68597a0ffffe780207e00005a85d285cdbf5685a685f5b72685ddb72285ddbf5d7186e4a2e026fc8505a5c12a8408659314150063e39500ae84914563e39500914497b5000083b5a5e8b3b5b400930640063386d402860509c918603305d5023af0894636f42af811a002f42800141097b0ffffe780e0a5a265426581cdfd55fe158505630ab50009ed9750ffffe780402c000008e004e4a6600664e2746161828062659750ffffe780002a0000130101dc233c1122233881222334912223302123233c312123384121368483c60600ba84b2892e8a2a89e5ce83c5040085e11385140097f5feff9385a5df1306000297a00000e78020b50125630905140a8597200000e78060ad0545230ca1100a852c0a05469760ffffe780e0aa230c41110a852c0a05469760ffffe780c0a90a8513060002ce859760ffffe780c0a8280aa28597000000e78080130a852c0a130600029760ffffe78000a7280aa68597000000e780c0110a852c0a130600029760ffffe78040a5280a8a851306800f97900000e780c0691304190002ea02e602e282fd280aac199770ffffe780605fac1913060002228597900000e7804067230009008330812303340123833481220339012283398121033a01211301012482801305140097f5feff9385a5d01306000297a00000e78020a683c5040001253366b50029e61385140097f5feff938565ce1306000297a00000e780e0a301250de9130610024a8581458330812303340123833481220339012283398121033a0121130101241793000067008351e31105ea05474a85d2854e86a68631a04a85d2854e86a28601478330812303340123833481220339012283398121033a012113010124170300006700e30f130101dc233c1122233881222334912223302123233c3121ae8483c505002a89d5c51384240093892402280097200000e780009309452300a11228000c1205469760ffffe7808090280013060002a2859760ffffe780808f280013060002ce859760ffffe780808e038514002300a11228000c1205469760ffffe780208d08122c001306800f97900000e780a05102ee02ea02e602e208120c029770ffffe78080470c02130600024a8597900000e780604f833081230334012383348122033901228339812113010124828093851400130600024a85833081230334012383348122033901228339812113010124179300006700234b130101da233c1124233881242334912423302125233c312323384123b68483c606002e892a84638a061403c5b40383c5a40303c6c40383c6d40322054d8d4206e206558e518d83c5f40303c6e40383c6040483c71404a205d18dc206e207dd8ed58d82154d8daaea03c5340383c5240303c6440383c6540322054d8d4206e206558e518d83c5740303c6640383c6840383c79403a205d18dc206e207dd8ed58d82154d8daae603c5b40283c5a40203c6c40283c6d40222054d8d4206e206558e518d83c5f40203c6e40283c6040383c71403a205d18dc206e207dd8ed58d82154d8daae203c5340283c5240203c6440283c6540222054d8d4206e20683c57402558e518d03c66402a20583c6840283c794024d8e93852400c206e207dd8e558e0216518d2afe05c3131589036d91301a329503060500937679000547b316d700558e2300c500130524001306000297900000e780c035130524022c1a1306000297900000e780a034038514000525a300a40005452300a4007da8b289850402ec02e802e402e005c3131589036d918a852e95830505001376790085463396c600d18d2300b500130a2400081097100000e780a06b230c211308102c1a054605499750ffffe7802069081013060002ce859750ffffe7802068081013060002a6859750ffffe7802067281a0c101306800f97900000e780a02b02fa02f602f202ee281a2c0a9770ffffe78080212c0a13060002528597900000e7806029130524028a851306000297900000e7804028a3002401230024018330812503340125833481240339012483398123033a0123130101268280157186eda2e9a6e5cae14efd52f956f55af15eed62e966e5328a7d16637ab63c2e89637aba3aaa89930a7102130b7108930b7108130c71065284050a93146400ce9403c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8d2ae103c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8daafc03c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8daaf803c5140083c5040003c6240083c6340022054d8d4206e206558e518d83c5540003c6440083c6640003c77400a205d18dc2066207d98ed58d82154d8daaf403c594fd83c584fd03c6a4fd83c6b4fd22054d8d4206e206558e518d83c5d4fd03c6c4fd83c6e4fd03c7f4fda205d18dc2066207d98ed58d82154d8d2af003c514fd83c504fd03c624fd83c634fd22054d8d4206e206558e518d83c554fd03c644fd83c664fd03c774fda205d18dc2066207d98ed58d82154d8d2aec03c594fc83c584fc03c6a4fc83c6b4fc22054d8d4206e206558e518d83c5d4fc03c6c4fc83c6e4fc03c7f4fca205d18dc2066207d98ed58d82154d8d2ae803c514fc83c504fc03c624fc83c634fc22054d8d4206e20683c554fc558e518d03c644fca20583c664fc03c774fcd18d938c04fcc2066207d98ed58d82154d8d2ae40155da855686630b051883c60500034706007d16fd150505e387e6fe63f0e618280013060004a68597900000e78080ff130600042685e68597900000e78080fe7d14630504147d1493146400ce940275e2654266a266aaf0aeecb2e8b6e403c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8d2ae103c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8daafc03c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8daaf803c5140083c5040003c6240083c6340022054d8d4206e206558e518d83c5540003c6440083c6640003c77400a205d18dc2066207d98ed58d82154d8daaf40155e2855e8605c983c60500034706007d16fd150505e388e6fe63fee600130600046685a68597900000e78040eaa68ce31004ecce8c2c0013060004668597900000e780c0e8e3132ac7ee604e64ae640e69ea794a7aaa7a0a7bea6b4a6caa6c2d61828017e5feff130585599305e0029790ffffe78000580000317106fd22f926f54af14eed52e956e55ae1defce2f8e6f4eaf02e89aa8993da1500130bf103930bf101130cf103930cf101fd1a13961a00130816006377284956850906637f262193166800ce9603c7960183c7860183c4a60103c4b60122075d8fc2046204458c418f83c7d60183c4c60103c4e60183c5f601a207c58f4204e205c18ddd8d8215d98d2eec83c5160103c7060183c7260183c43601a205d98dc207e204c58fdd8d03c7560183c7460183c4660103c4760122075d8fc2046204458c418f0217d98d2ee883c5960003c7860083c7a60083c4b600a205d98dc207e20403c7d60003c4c600c58fdd8d2207418f83c7e60083c4f6001a064e96c207e204c58f5d8f0217d98d2ee483c5160003c7060083c7260083c43600a205d98dc207e204c58fdd8d03c7560083c7460083c4660083c6760022075d8fc204e206c58ed98e8216d58d2ee083459601834686010347a6018347b601a205d58d4207e2075d8fd98d8346d6010347c6018347e6018344f601a206d98ec207e204c58fdd8e8216d58d2efc83451601834606010347260183473601a205d58d4207e2075d8fd98d83465601034746018347660183447601a206d98ec207e204c58fdd8e8216d58d2ef883459600834686000347a6008347b600a205d58d4207e2075d8fd98d8346d6000347c6008347e6008344f600a206d98ec207e204c58fdd8e8216d58d2ef483451600834606000347260083473600a205d58d4207e2075d8fd98d83465600034746008347660003467600a206d98ec20762065d8e558e0216d18d2ef00156de865a8719ce83c70600834407007d17fd160506e38897fe33ba970021a0428a19a0014a429a6379257763742a771a053384a90093146a00ce9403459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8d2aec0345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8d2ae803459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8d2ae40345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8d2ae003c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8d2afc03c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8d2af803c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8d2af403c5140083c5040003c6240083c6340022054d8d4206e206558e518d83c5540003c6440083c6640003c77400a205d18dc2066207d98ed58d82154d8d2af00155e685628639c983c60500034706007d16fd150505e388e6fe63f1e604081013060004a28597900000e780c09b130600042285a68597900000e780a0df0c1013060004268597900000e780c09913161a00130816005285e36e28b7e3940ab6130bf103930bf101130cf103930cf101094dca8afd1a63fb2a4f13946a004e94081013060004ce8597900000e780a095130600044e85a28597900000e78080d90c1013060004228597900000e780a09363ebaa490146014505480906637f562193166800ce9603c7960183c7860183c4a60103c4b60122075d8fc2046204458c418f83c7d60183c4c60103c4e60183c5f601a207c58f4204e205c18ddd8d8215d98d2eec83c5160103c7060183c7260183c43601a205d98dc207e204c58fdd8d03c7560183c7460183c4660103c4760122075d8fc2046204458c418f0217d98d2ee883c5960003c7860083c7a60083c4b600a205d98dc207e20403c7d60003c4c600c58fdd8d2207418f83c7e60083c4f6001a064e96c207e204c58f5d8f0217d98d2ee483c5160003c7060083c7260083c43600a205d98dc207e204c58fdd8d03c7560083c7460083c4660083c6760022075d8fc204e206c58ed98e8216d58d2ee083459601834686010347a6018347b601a205d58d4207e2075d8fd98d8346d6010347c6018347e6018344f601a206d98ec207e204c58fdd8e8216d58d2efc83451601834606010347260183473601a205d58d4207e2075d8fd98d83465601034746018347660183447601a206d98ec207e204c58fdd8e8216d58d2ef883459600834686000347a6008347b600a205d58d4207e2075d8fd98d8346d6000347c6008347e6008344f600a206d98ec207e204c58fdd8e8216d58d2ef483451600834606000347260083473600a205d58d4207e2075d8fd98d83465600034746008347660003467600a206d98ec20762065d8e558e0216d18d2ef00156de865a8719ce83c70600834407007d17fd160506e38897fe33ba970021a0428a19a0014a429a63715529637e5a271a053384a90093146a00ce9403459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8d2aec0345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8d2ae803459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8d2ae40345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8d2ae003c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8d2afc03c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8d2af803c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8d2af403c5140083c5040003c6240083c6340022054d8d4206e206558e518d83c5540003c6440083c6640003c77400a205d18dc2066207d98ed58d82154d8d2af00155e6856286e30405b883c60500034706007d16fd150505e387e6fee3f9e6b6081013060004a28597800000e780404d130600042285a68597900000e78020910c1013060004268597800000e780404b13161a00130816005285e36d58b705beea704a74aa740a79ea694a6aaa6a0a6be67b467ca67c067d296182805285d68529a0528511a05685ca859790ffffe780c0430000757106e522e1a6fccaf8cef4d2f0d6ecdae8dee4ae89fd1513d61500d18d13d62500d18d13d64500d18d13d68500d18d13d60501d18d13d60502d18d93c5f5ff17a60000033626ae97a6000083b626ae13d71500798e918d33f6d5008981f58db29517a60000033606ad97a6000083b606ad13d74500ba95f18db385d502e1917d56b35ab600850a638a0a0a2a8913d519007999fd1a130bf5ff13d529001e054a95130405fc8d44ce8b63723b091395db0033457501935575002d8d93151501b3cba50033f55b01b3353501fd15b3f535010d8d637e35051a05330aa900280013060004a28597800000e7802038130600042285d28597800000e780007c2c0013060004528597800000e7802036050bfd1413040404d1f8aa600a64e6744679a679067ae66a466ba66b496182805a85ce859790ffffe7800030000017e5feff1305e5a3f1459790ffffe78080a40000557186e5a2e126fd4af94ef552f156ed5ae95ee562e1e6fceaf8eef42e8c2a89014b930b7104930c710213bd2503954d854463f384238545139564004a9503469501834685010347a5018347b5012206558e4207e2075d8f598e8346d5010347c5018347e5010344f501a206d98ec2076204c18fdd8e8216558e32f0034615018346050103472501834735012206558e4207e2075d8f598e83465501034745018347650103447501a206d98ec2076204c18fdd8e8216558e32ec03469500834685000347a5008347b5002206558e4207e2075d8f598e8346d5000347c5008347e5000344f500a206d98ec2076204c18fdd8e8216558e32e8034615008346050003472500834735002206558e4207e2075d8f598e83465500034745008347650003447500a206d98ec2076204c18fdd8e8216558e32e4034695fd834685fd0347a5fd8347b5fd2206558e4207e2075d8f598e8346d5fd0347c5fd8347e5fd0344f5fda206d98ec2076204c18fdd8e8216558eb2e0034615fd834605fd034725fd834735fd2206558e4207e2075d8f598e834655fd034745fd834765fd034475fda206d98ec2076204c18fdd8e8216558e32fc034695fc834685fc0347a5fc8347b5fc2206558e4207e2075d8f598e8346d5fc0347c5fc8347e5fc0344f5fca206d98ec2076204c18fdd8e8216558e32f8034615fc834605fc034725fc834735fc2206558e4207e2075d8f598e834655fc034745fc834765fc034575fca206d98ec20762055d8d558d0215518d2af401556686de8601cd0347060083c70600fd167d160505e308f7fe6369f7008504b3b58401e39384df51a0814533c58401133515003366ad003dea9389f4ff63f789098589d1c5139a69004a9a939a6400ca9a281013060004d28597800000e7800009130600045285d68597800000e78000082c1013060004568597800000e78000070545637f95004a85a6854e8697f0ffffe78060e04a85a68597000000e7804004050be310bbd7014511a00545ae600e64ea744a79aa790a7aea6a4a6baa6b0a6ce67c467da67d696182804e8511a02685e2859790ffffe78000fe0000317106fd22f926f54af14eed52e956e55ae12e89aa840345950583c5840503c6a40583c6b40522054d8d4206e206558e518d83c5d40503c6c40583c6e40503c7f405a205d18dc2066207d98ed58d82154d8daafc03c5140583c5040503c6240583c6340522054d8d4206e206558e518d83c5540503c6440583c6640503c77405a205d18dc2066207d98ed58d82154d8daaf803c5940483c5840403c6a40483c6b40422054d8d4206e206558e518d83c5d40403c6c40483c6e40403c7f404a205d18dc2066207d98ed58d82154d8daaf403c5140483c5040403c6240483c6340422054d8d4206e206558e518d83c5540403c6440483c6640403c77404a205d18dc2066207d98ed58d82154d8daaf003c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8d2aec03c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8d2ae803c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8d2ae403c5140083c5040003c6240083c6340022054d8d4206e20683c55400558e518d03c64400a20583c6640003c77400d18d93890404c2066207d98ed58d82154d8d2ae01305f10181551306f1076380051a83460600034705007d157d168505e387e6fe63f5e6180a8513060004a68597800000e78060dd130600042685ce8597800000e78060dc0d45636aa914130af107894a130bf10513946a00269403459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8daaec0345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8daae803459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8daae40345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8daae06265c26522668266aafcaef8b2f4b6f00155da8552860dc983c60500034706007d16fd150505e388e6fe63ffe600850a130504fc13060004a28597800000e78060c7a289e39f2aeb8a85130600044e8597800000e78000c6ea704a74aa740a79ea694a6aaa6a0a6b29618280257106ef22eb26e74ae32a8484004800130901031306c002814597800000e780c0b5130680132685814597800000e780c0b417d5feff9305550741464a8597800000e78060c0370501011b0505022ac082fe8a8522859740ffffe78000e4fa605a64ba641a691d6182805d7186e4a2e026fc8505a5c12a8408659314150063e39500ae84914563e3950091449795000083b52529b3b5b400930600053386d4028e0509c918603305d5023af0a14636f42af811a002f4280014109790ffffe780e0e3a265426581cdfd55fe158505630ab50009ed9730ffffe780406a000008e004e4a6600664e2746161828062659730ffffe780006800005d7186e4a2e026fc4af8ae84806590612a892800a2859770ffffe78080400345810001c9426505c59780ffffe7806041000005040dc49305910080e4130519001306000297800000e78080b005452300a900a6600664e27442796161828017d5feff13050520f1459780ffffe780a02000000e0597d5feff938525962e950c6105458285094582800d458280114582809780ffffe780e03a0000106195456316b60003058500050582800c65328517030000670043fc130101d32334112c2330812c233c912a2338212b2334312b2330412bb2842e842a8902f002ec02e802e4930901164812130a01151306c002814597800000e780e098130680134e85814597800000e780e09717d5feff930575ea4146528597800000e78080a3370501011b0505022320a112233c012828100c129740ffffe780e0c62810a28526869740ffffe78060db08122c101306800f97800000e780e09f08122c009760ffffe78040962c00130600024a8597800000e780209e8330812c0334012c8334812b0339012b8339812a033a012a1301012d8280317106fd22f926f54af14eed52e993070002631cf61eba89368a2a8903c5950103c6850183c6a50103c7b5012205518dc2066207d98e558d03c6d50183c6c50103c7e50183c7f5012206558e4207e2075d8f598e0216518d2aec03c5150103c6050183c6250103c735012205518dc2066207d98e558d03c6550183c6450103c7650183c775012206558e4207e2075d8f598e0216518d2ae803c5950003c6850083c6a50003c7b5002205518dc2066207d98e558d03c6d50083c6c50003c7e50083c7f5002206558e4207e2075d8f598e0216518d2ae403c5150003c6050083c6250003c735002205518dc2066207d98e558d03c6550083c6450003c7650083c575002206558e4207e205d98dd18d82154d8d2ae088009770ffffe78040c6a8188a859770ffffe78000b3266511c506659730ffffe780e0392a658a6566762afc2ef832f40305710783056107e664034651072303a102a20503452107d18d2312b10283451107220503463107830641074d8d06744206e206558e518d2ad0a818d2854e869770ffffe780e0b111c426859730ffffe780e0332275e6754276aae062758a66b2e42a66aae8aeecb6f0b2f405452308a106130511070c101d4697700000e780e07fa8188c009770ffffe78020c3880097000000e780600566742a664a85a28597000000e78020d40a6511c522859730ffffe780c02dea704a74aa740a79ea694a6a2961828017d5feff130525f197d5feff9386c5f39305b00290009780ffffe78020070000411106e422e02a84086511c508609730ffffe7806029087009c9086ca260026441011733ffff67002328a260026441018280697106f622f226ee4aea4ee652e2d6fddaf9def5e2f1e6ed2e8a2a89014481490d45aae082e49304110501163335c00093b51500b36ab500130b1108894b7d5c88088c009790ffffe780a051034501056309751f6301051003c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8d2ae903c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8d2ae503c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8d2ae103c5140083c5040003c6240083c6340022054d8d4206e206558e518d83c5540003c6440083c6640003c77400a205d18dc2066207d98ed58d82154d8daafc63890a00dda002e902e502e182fc639e0a0ca81813060002d28597800000e780e0a1012579e1639a091628110d46a2859770ffffe780e0fa2a7559c96a75ca752a76aae9aee5b2e1a8188c019790ffffe78020220305eb008305db000346cb00e6792303a10aa205d18d2312b10a03459b0083458b000346ab008306bb0022054d8d4206e206558e518d2ad103451b0083450b0003462b0083463b0022054d8d4206e20683455b00558e518d03464b00a20583466b0003477b00d18d834c0108c2066207d98ed58d82154d8d2aed11a081496a658a550316410a8306610a2af82edc231ec102230fd102630e8409050401b5638609060305e1038315c1036256c2762307a1022316b10232d436f0130511010c103d4697700000e780a04f4ee423089101a8182c0005469790ffffe78080d6667535c92a658a656676aaf0aeecb2e888089790ffffe78080f12334a9004e859790ffffe78060a4014531a01305a005a300a90005452300a900b2701274f2645269b269126aee7a4e7bae7b0e7cee6c5561828017d5feff1305c5b9f1459780ffffe78060ba000017d5feff130585ec9305b002edb717d5feff130585bc97c5feff9386253c9305b00290089780ffffe78080d20000497186f6a2f2a6eecaeacee6d2e256fe5afa5ef662f266ee6aea6ee62e842ae0814a014d0149014b0945aaf882fc93041108bd497d5a2ee408018c1897000000e780008c03450108630b052803c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8daae103c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8d2afd03c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8d2af903c5140083c5040003c6240083c6340022054d8d4206e206558e518d83c5540003c6440083c6640003c77400a205d18dc2066207d98ed58d82154d8d2af5281113060002a28597700000e780407201256310051888190946d6859770ffffe78060cbce7b638a0b1e126c6e7563fc8915aae8eaec414581459780ffffe78060642a842e8b4146de8597700000e780a02b83458400834994000349a400834db4000346c400034dd4008347e400034af400834c04000347140083432400834634000348440003435400834864008342740063050b04228542f0468416fc6aec1a8d4ae81e896ef4b68dcee0ba89b2e452f83e8a2e8b9730ffffe78000d6da85d287427a26664e878669ee86a27dca8342696a83626de272a28802786665631e0514a20933e5b9004209e20db3e52d014d8d220db365cd0013960701620a3366ca00d18d8215b3eda50013158700336595019395030113968601d18d4d8d93158300b3e505011396080193968201558ed18d8215b3eca50013040cff93890b01228581459780ffffe780c0532a8c2e8bce85228697700000e780001be2f9dafd22e2a8098c199790ffffe780c0df8c1188618c65014b6e6daaf0aef405492264bd497d5a466511c55e859730ffffe780c0c8638a4a07850ab1bb3365690119cd630d0d0226758675026608f20cee233096012334b6012338a6013da01305500382652380a50023b80500630f0d006a859780ffffe780c06b01a81305200382652380a50023b80500b6701674f6645669b669166af27a527bb27b127cf26c526db26d7561828017d5feff13050581f1459780ffffe780a081000017d5feff1305a58497d5feff938645899305b002b0099780ffffe780a09a000017d5feff130575b493059002e9b7097186fea2faa6f6caf2ceeed2ead6e6dae25efe62fa66f66af26eeeb289ae842ae4014b014d0149814b32e102e5130411093d4afd5a32ec2ee808090c0197f0ffffe780205303450109630c052803459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8daae90345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8daae503459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8daae10345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8d2afd281913060002a68597700000e78060390125631105180802da854e869770ffffe7808092126c630b0c1ed26c3265637d9a15aaf0eaf4414581459780ffffe780802baa84ae8b4146e28597700000e780c0f283c5840003ca940003c9a40083c9b40003c6c40083cdd40083c7e40083caf40003cd040003c7140083c3240083c6340003c8440003c3540083c8640083c2740063850b042685c28bc684d6e016f86ef49a8d4af01e89b6e4d2e83a8ab2ec4efcbe89ae8a9730ffffe780209dd685ce87e27966665287466aa666ca8302796e83a27dc272866aa6885e882675631f0514220a3365ba004209e209b3e529014d8da20db3e5cd0013960701e20a33e6ca00d18d82154d8daaf4131587003365a5019395030113968601d18d4d8d93158300b3e505011396080193968201558ed18d8215b3eda50093840cff130a0c01268581459780ffffe780e01aaa8cae8bd285268697700000e78020e266e25ee626eaa8110c029790ffffe780e0a68c1988618c65814b2e7daaf8aefc0549e269c2643d4afd5a067511c562859730ffffe780c08f630a5b07050ba9bb3365790119cd630d0d026675c675226608f20cee2330b601267508e62338a6013da013055003a2652380a50023b80500630f0d006a859780ffffe780c03201a813052003a2652380a50023b80500f6705674b6741679f669566ab66a166bf27b527cb27c127df26d1961828017c5feff13050548f1459770ffffe780a048000017c5feff1305a54b97c5feff938645509305b002b0119770ffffe780a061000017c5feff1305057e9305c002e9b7097186fea2faa6f6caf2ceeed2ead6e6dae25efe62fa66f66af26eeeae892ae4014b814a214a52e802ec02f005452af402f8130d9103930d110b0944fd5428182c109790ffffe78080ae034581036309853475cd03459d0183458d010346ad018346bd0122054d8d4206e206558e518d8345dd010346cd018346ed010347fd01a205d18dc2066207d98ed58d82154d8daae503451d0183450d0103462d0183463d0122054d8d4206e206558e518d83455d0103464d0183466d0103477d01a205d18dc2066207d98ed58d82154d8daae103459d0083458d000346ad008346bd0022054d8d4206e206558e518d8345dd000346cd008346ed000347fd00a205d18dc2066207d98ed58d82154d8d2afd03451d0083450d0003462d0083463d0022054d8d4206e206558e518d83455d0003464d0083466d0003477d00a205d18dc2066207d98ed58d82154d8d2af929a082e582e102fd02f9081913060002ce8597700000e78060ff01256318052208190546da859760ffffe780c0480345010b6311052603c59d0183c58d0103c6ad0183c6bd0122054d8d4206e206558e518d83c5dd0103c6cd0183c6ed0103c7fd01a205d18dc2066207d98ed58d82154d8daafc03c51d0183c50d0103c62d0183c63d0122054d8d4206e206558e518d83c55d0103c64d0183c66d0103c77d01a205d18dc2066207d98ed58d82154d8daaf803c59d0083c58d0003c6ad0083c6bd0022054d8d4206e206558e518d83c5dd0003c6cd0083c6ed0003c7fd00a205d18dc2066207d98ed58d82154d8daaf403c51d0083c50d0003c62d0083c63d0022054d8d4206e206558e518d83c55d0003c64d0083c66d0003c77d00a205d18dc2066207d98ed58d82154d8daaf008190546da859760ffffe780a047ca7b63870b168e653d456378b51a6a79138405ff138c0b01228581459780ffffe78040e0aa84ae8ce285228697700000e78080a726f966fda2e108010c199780ffffe780406c28090c019730ffffe780609608020c010d469780ffffe780e02c1265630305125265b2651266aae12efd32f908020c199780ffffe78000575265d145631cb510126451468809a28597700000e78060a13265fd5411c522859720ffffe78080510675a67546762af92efdb2e16675aa750a76ea666267aae5a8110ce910e514e1639aea000808d68597f0ffffe780c0df827a426a0944130500053385aa0252950c191306000597700000e780809b0a65850a56f09780ffffe78020f3630709005e859720ffffe780e04a630a9b02050b45b10275e2654266a26688ea8ce690e2f6705674b6741679f669566ab66a166bf27b527cb27c127df26d1961828017c5feff13052507f1459770ffffe780c007000017c5feff1305c50a97c5feff9386650f9305b002901089a017c5feff1305450997c5feff9386e50d9305b00210022da017c5feff1305c50797c5feff9386658709a817c5feff1305a50697c5feff938645099305b00210199770ffffe780a01c000041459780ffffe780208b0000757106e522e1a6fccaf8cef4d2f02a89814432e402e81304910181153335b00093351900b369b500094a28082c009780ffffe780e06a0345810165d9630c451303459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8daaec0345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8daae803459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8daae40345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8daae0e39909ee880013060002ca8597700000e78020bc0125e31e05ec93f4f40f850413f5f40fe30795ec17c5feff130505e9f1459770ffffe780a0e900002685aa600a64e6744679a679067a49618280517186f5a2f1a6edcae9cee5d2e156fd5af95ef562f166ed6ae96ee5b2892e8a2ae0014b814a32ec02f013049102894d7d5928102c089780ffffe7800052034581026300b51b75cd03459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8daaf40345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8daaf003459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8daaec0345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8daae829a082f482f082ec82e8880813060002d28597700000e780e0a2012519c1d684a5a88808da854e869760ffffe780e0fbc66b63820b0c666d8674268581459780ffffe7806095aa8c2e8cde85268697600000e780a05ce6e8e2eca6f088188c089780ffffe7806021ac1888618c65c674aae8aeec63870a0056859780ffffe78060b26665c6652ae82ee463070d005e859720ffffe780a00963052b05050ba68a89bd63890a004265a265026608ea32850ce639a01305b00682652384a5002e8523305501ae700e74ee644e69ae690e6aea7a4a7baa7b0a7cea6c4a6daa6d6d61828017c5feff130585c4f1459770ffffe78020c5000017c5feff130525c897c5feff9386c5cc9305b00290189770ffffe78020de00001d7186eca2e8a6e4cae02a84081097000000e780c0d98274a1c40309810293059102130511013d4697600000e780a04d26e42308210108102c000d469780ffffe78080d402750dc94275a275027608e80ce410e026859780ffffe78040a339a0030581022304a40023300400e6604664a66406692561828017c5feff1305a5be97b5feff9386453e9305b0021306f1039770ffffe78080d40000357106ed22e926e5aa85a8100d4697000000e78020d0267461c88304010793051107130511013d4697600000e780004422e423089100a8102c0011469780ffffe780e0ca26754dcd6675c67526762af82ef432f0a8100c1001469780ffffe78000c926755dc56675c6752676aae4aee032fc88082c1809469780ffffe78020c7466545c50675e6654666aafcaef8b2f4231201088808ac105001894689449780ffffe780809a0345010541ed6665631b950a8314410826759780ffffe780809362759780ffffe780e09202759780ffffe780409222859780ffffe780a091014501469b95040131a003450107814522050546d18d4d8dea604a64aa640d61828017c5feff130585ac97b5feff9386252c09a817c5feff130565ab97b5feff9386052b9305b00290080da817c5feff1305e5a997b5feff938685299305b002b01029a817c5feff130565a897c5feff938605809305b002130671089770ffffe78040be000017c5feff1305c591b9459770ffffe78000a20000517186f5a2f1a6edcae9cee5d2e156fd5af95ef562f166ed6ae96ee5b2892e8a2ae0014b814a32ec02f013049102894d7d5928102c089780ffffe780800b034581026300b51b75cd03459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8daaf40345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8daaf003459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8daaec0345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8daae829a082f482f082ec82e8880813060002d28597600000e780605c012519c1d684a5a88808da854e869760ffffe78060b5c66b638a0b0a666d8674268581459770ffffe780e04eaa8c2e8cde85268697600000e7802016e6e8e2eca6f088188c089780ffffe780e0daac1888618c65c674aae8aeec63870a0056859770ffffe780e06b6665c6652ae82ee463070d005e859720ffffe78020c3630d2b03050ba68a89bd63820a064265a265026608ea0ce623305601ae700e74ee644e69ae690e6aea7a4a7baa7b0a7cea6c4a6daa6d6d61828017b5feff1305057ff1459760ffffe780a07f000017c5feff1305a58297c5feff938645879305b00290189770ffffe780a098000017b5feff1305e5789305b002e9b7130101ce233c1130233881302334913023302131233c312f2338412f2334512f2330612f233c712d2338812d2334912d2330a12d233cb12b3a8a3684328bae892a891305000285459720ffffe780e0b56306056eaa8413060002814597600000e78020f7514585459720ffffe780e0b36309056c2a8c5146814597600000e78040f51305000281459770ffffe7800039aa8bae8a13060002d28597600000e780200026859720ffffe780a0b00345140183450401034624018306340122054d8d4206e206558e518daac803459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8daae40345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8daae0130a0105930c8104514581459770ffffe780602c2afeaee282e693041104281a8c0026869770ffffe780601113042104281aa68522869770ffffe780401093043104281aa28526869770ffffe780200fc000281aa68522869770ffffe780200e93045104281aa28526869770ffffe780000d13046104281aa68522869770ffffe780e00b93047104281aa28526869770ffffe780c00a281aa68566869770ffffe780e00913049104281ae68522869770ffffe780c0089304a104281aa28526869770ffffe780a0071304b104281aa68522869770ffffe7808006e400281aa28526869770ffffe78080051304d104281aa68522869770ffffe78060049304e104281aa28526869770ffffe78040031304f104281aa68522869770ffffe7802002281aa28552869770ffffe780400113041105281ad28522869770ffffe780200093042105281aa28526869770ffffe78000ff13043105281aa68522869770ffffe780e0fdd008281aa2859770ffffe78000fdf27c966d366a62859720ffffe780e08e1304ca02636e4445228581459770ffffe78040142afeaee282e64145a1459720ffffe780008c630c05442a8c31452330ac001305c0022334ac00a2c0d000281a8c009770ffffe78060f78944130d410462840860aac0281a8c006a869770ffffe780c0f5fd142104edf462859720ffffe780a08713860b02281ade859770ffffe780c0f333864c01281ae6859770ffffe780c0f2727a166d366c63870a005e859720ffffe780608463870d0066859720ffffe78080835a8581459770ffffe78060092a84ae8ace855a8697600000e780a0d013050002631aab3a03056400230fa112030554008345440022054d8d231ea1120345140083450400034624008306340022054d8d4206e206558e518d232ca1120345840083457400034694008346a40022054d8d4206e206558e518d8345c4000346b4008346d4000347e400a205d18dc2066207d98ed58d8215b3e9a500034504018345f400034614018346240122054d8d4206e206558e518d83454401034634018346540103476401a205d18dc2066207d98ed58d8215b3eba5000345840183457401034694018346a40122054d8d4206e206558e518d8345c4010346b4018346d4010347e401a205d18dc2066207d98e034bf401d58d8215b3e4a50063870a0022859710ffffe78000710305e1138315c113032681132303a1042312b104b2c0a303310513d589032307a10413d50903a306a10413d589022306a10413d50902a305a10413d589012305a10413d50901a304a10413d589002304a104a307710513d58b03230ba10413d50b03a30aa10413d58b02230aa10413d50b02a309a10413d58b012309a10413d50b01a308a10413d58b002308a104a30b910413d58403230fa10413d50403a30ea10413d58402230ea10413d50402a30da10413d58401230da10413d50401a30ca104a180230c9104a30f6105281a9750ffffe78060ee08108c009750ffffe78020db166511c572759710ffffe78000624275a27502762aec2ee832e40305f1168305e11656640346d1162303a100a2050345a116d18d2312b1008345911622050346b1168306c1164d8df6644206e206558e518d2ac00810d28562869750ffffe78000da91c422859710ffffe780005c2265827542662afe6265a276b2e24276aae6aeeab6eeb2f205452304a116130591168a851d4697600000e78000a828002c1a9750ffffe78040eb281a97e0ffffe780802d02fc02f802f402f0a01a681aa4121306c002814597600000e7800098130680132285814597600000e780009717b5feff930595e94146268597600000e780a0a2370501011b050502232ca1122338012a88002c1a9720ffffe78000c6226462668800a2859720ffffe78060da281a8c001306800f97600000e780e09e281a0c109740ffffe78040950c10130600024a8597600000e780209d426511c522859710ffffe780604d63070d0052859710ffffe780804c833081310334013183348130033901308339812f033a012f833a812e033b012e833b812d033c012d833c812c033d012c833d812b13010132828017b5feff1305658ff1459760ffffe780000900001305000221a0514511a041459710ffffe780e047000017b5feff1305a50a97b5feff938645119305b002301a9760ffffe780a0200000130101dd2334112223308122233c91202e84aa8402f002ec02e802e4281097e0ffffe78080cc22f228100c1221469720ffffe78040ca08122c101306800f97600000e780c08e08122c009740ffffe78020852c0013060002268597600000e780008d833081220334012283348121130101238280130101812334117e2330817e233c917c2338217d2334317d2330417d233c517b2338617b2334717b2330817b233c91792338a1792334b179357136ec32e42ee82a842338014623340146a80813068002814597500000e78060790335014683358146033601472ae12ee5086032e902f10c683336a00014643307c040f98d32f502f92afdb6e1b2e582e9aaedb6f1aef5130da122930ba124854d930a400828119770ffffe780606819e16f2090222a8493040501233c0178233801782334017823300178881697e0ffffe780c0ba88165146a6859720ffffe780a0b8130501468c161306800f97500000e780007d13050146930501789730ffffe7802073033581798335017903368178833601782ae62ee2b2fdb6f9033b0400033c84002af62ef232ee36ea233c0178233801782334017823300178881697e0ffffe780a0b3233481472330614788169305014641469720ffffe780e0b0130501468c161306800f97500000e780407513050146930501789730ffffe780606b930501781306000213041113228597500000e780e0722308011217b5feff930565de13060002228597600000e780c0b3012521c1327592757266d2664a6a2334a1282330b128233cc1262338d12663080a046a648c1c52859770ffffe7808077ae842dcd41c48e04d29403ba04227d14d5b74a64e30a04386a65b384ad400c0a22859770ffffe780e07463000518e38db4378e05a29503b405228504cdb7833981278334012803398128033401279770ffffe780e05b233805208545231db52000e12334350104e9233c250123348517233065172ae902ed6f00f0329204d29423b4841723b064176f001032033d812783350128833c81280359aa21833b01272d456379a91293891400139454005294939a44006375391d2300740113d58b03a303a40013d50b032303a40013d58b02a302a40013d50b022302a40013d58b01a301a40013d50b012301a40013d58b00a300a4002304a40113558d03a307a40013550d032307a40013558d02a306a40013550d022306a40013558d01a305a40013550d012305a40013558d00a304a4002308b40013d58503a30ba40013d50503230ba40013d58502a30aa40013d50502230aa40013d58501a309a40013d505012309a40013d58500a308a400230c940113d58c03a30fa40013d50c03230fa40013d58c02a30ea40013d50c02230ea40013d58c01a30da40013d50c01230da40013d58c00a30ca400f5aa2300015a639ab40323308136233401362338b136130501468c161306015a9770ffffe78040616f20206f854d1545aee463f2a41e1149e5aa8e05a29503b5052299c8b30590400356a5210e06329503350522fd15edf98355a521fd152338a164233c01642330b16613050146930501651306015a9770ffffe780e05b0335814783350147233ca17803368146833601462338b178033501492334c1782330d1780339014a8355a521833481492a846374b9006f20004e0334052119e06f20204d035985218355a42185042285e375b9fe6f20204c139559005295b304994013965400d6e8ae8aa28597600000e780808913d58b03a303a40013d50b032303a40013d58b02a302a40013d50b022302a40013d58b01a301a40013d50b012301a40013d58b00a300a4002300740113558d03a307a40013550d032307a40013558d02a306a40013550d022306a40013558d01a305a40013550d012305a40013558d00a304a4002304a40113d58a03a30ba40013d50a03230ba40013d58a02a30aa40013d50a02230aa40013d58a01a309a40013d50a012309a40013d58a00a308a40023085401c66a13d58c03a30fa40013d50c03230fa40013d58c02a30ea40013d50c02230ea40013d58c01a30da40013d50c01230da40013d58c00a30ca400230c940113050a16b305550192094e951396440097500000e780e0780529d29a23b48a1723b06a17231d2a21130da122930ba124cda76389a400814d19456397a4008144154929a0268919a0e5141949e2e09770ffffe7802023aa8a23380520231d05200355aa219349f9ffaa99239d3a2193155900d29503c6950183c6850103c7a50183c7b5012206558e4207e2075d8f598e83c6d50103c7c50183c7e50103c4f501a206d98ec2076204c18fdd8e8216558e233cc14603c6150183c6050103c7250183c735012206558e4207e2075d8f598e83c6550103c7450183c7650103c47501a206d98ec2076204c18fdd8e8216558e2338c14603c6950083c6850003c7a50083c7b5002206558e4207e2075d8f598e83c6d50003c7c50083c7e50003c4f500a206d98ec2076204c18fdd8e8216558e2334c14603c6150083c6050003c7250083c735002206558e4207e2075d8f598e83c6550003c7450083c7650083c57500a206d98ec207e205dd8dd58d8215d18d2330b146b14563e4b9006f30802dca8613041900018d630435016f30e02c5a8c6689930c0a161395460066950c65aee808612afc93155400d295139659005685368b97500000e780e01993154400e69513850a161396490097500000e7808018231d6a21033501468335814603360147833681472330a1362334b1362338c136233cd136528663930d0056860357a6219389140013945400329493974400ca8c628b637c370f2300740113d58b03a303a40013d50b032303a40013d58b02a302a40013d50b022302a40013d58b01a301a40013d50b012301a40013d58b00a300a4002304a40113558d03a307a40013550d032307a40013558d02a306a40013550d022306a40013558d01a305a40013550d012305a40013558d00a304a400a6652308b40013d58503a30ba40013d50503230ba40013d58502a30aa40013d50502230aa40013d58501a309a40013d505012309a40013d58500a308a400230c940113d58c03a30fa40013d50c03230fa40013d58c02a30ea40013d50c02230ea40013d58c01a30da40013d50c01230da40013d58c00a30ca40005aa139559003295b30d9740328913965d00a2853a8cbe8497500000e780e04713d58b03a303a40013d50b032303a40013d58b02a302a40013d50b022302a40013d58b01a301a40013d50b012301a40013d58b00a300a4002300740113558d03a307a40013550d032307a40013558d02a306a40013550d022306a40013558d01a305a40013550d012305a40013558d00a304a4002304a401a66513d58503a30ba40013d50503230ba40013d58502a30aa40013d50502230aa40013d58501a309a40013d505012309a40013d58500a308a4002308b40013d58c03a30fa40013d50c03230fa40013d58c02a30ea40013d50c02230ea40013d58c01a30da40013d50c01230da40013d58c00a30ca400230c940113050916b305950092094e9513964d0097500000e7804037a68762874a86c66de27486661b051700b305f60023b4d51623b06517231da62003358137833501370336813683360136233ca1782338b1782334c1782330d178233ca15a2338b15a2334c15a2330d15a03350a216309052c8149d687268c6e8d03598a218335815b0336015b8336815a0337015a233cb1782338c1782334d1782a8a2330e178835ba5212d4563ebab32cee4054b91491545bee0636fa9006309a900014b19456317a9000149954929a0ca8919a0651999499770ffffe780e0dbaa8a23380520231d05200355aa2113c4f9ffb30ca400239d9a2193955900d29503c6950183c6850103c7a50183c7b5012206558e4207e2075d8f598e83c6d50103c7c50183c7e50183c4f501a206d98ec207e204c58fdd8e8216558e233cc14603c6150183c6050103c7250183c735012206558e4207e2075d8f598e83c6550103c7450183c7650183c47501a206d98ec207e204c58fdd8e8216558e2338c14603c6950083c6850003c7a50083c7b5002206558e4207e2075d8f598e83c6d50003c7c50083c7e50083c4f500a206d98ec207e204c58fdd8e8216558e2334c14603c6150083c6050003c7250083c735002206558e4207e2075d8f598e83c6550003c7450083c7650083c57500a206d98ec207e205dd8dd58d8215d18d2330b146b14563e4bc006f20505f93841900058d630495016f20d05e13040a161395490022950c65aee8833d050093955400d29513965c00568597500000e78080d093954400a29513850a1613964c0097500000e78020cf231d3a21033501462330a13603358146833501470336814783dcaa212334a1362338b136233cc13613851c00b14563e4bc006f20704c33863b416304a6006f209057a66985098e04d2949385042213840a220e06228597500000e78040c9014593153500a2958c6133369501239ca5203295b3b6ac0093c61600758e23b8552165f2033581378335013703368136833601362334a1662330b166233cc1642338d1645285866763130b00568513060178ca85e2866a879770ffffe78040bb033501658335816503360166833681662330a15a2334b15a2338c15a233cd15a03350a21d687ee846e8cc66d6e8de31005d411a081494a6419e06f2090516a699770ffffe78040b423380520231d052023308522930519002338a420231c04202ae92eed130da122930ba124630439016f20d04e8355a52129466374b6006f20904e1b861500231dc520139655008336015b2a960337015a8337815b14ea8336815a18e21cee1307052214e6139645002a96233096162334b6178505139635003a962330560123b8aa20239cba2039a8130601785285ca85e2866a879770ffffe78000ad130da122930ba124854d930a40088a7585052ef1327592757266d2662aeb2ee732e3b6fe280b0c1a1306200497500000e780c0b1034481177d461305111e9305911797500000e78060b0814c81491375e40f2300a11e05447e75de75233ca1203e751e762338b120667c2334a120a2e42330c120230031230949630a0c2a0a68e28283d8625b01451387825b93975800b30517013383f5001386725d63036706aa830345070293f5f90fb3b4a5002d8d3335a000b3059040c98d95e501541305f121b28421c88345050083c70400b3b6f500bd8db335b000b306d040d58dfd147d150504e5d1138513001307170213061602e385b5fb13f5f50f09cd631608003da4c683630508228e039e9283b282727d1885bf33855303169583458500930485006387052003c5b40183c5a40103c6c40183c6d40122054d8d4206e206558e518d83c5f40103c6e40183c6040203c71402a205d18dc2066207d98ed58d82154d8d233ca17803c5340183c5240103c6440183c6540122054d8d4206e206558e518d83c5740103c6640183c6840103c79401a205d18dc2066207d98ed58d82154d8d2338a17803c5b40083c5a40003c6c40083c6d40022054d8d4206e206558e518d83c5f40003c6e40083c6040103c71401a205d18dc2066207d98ed58d82154d8d2334a17803c5340083c5240003c6440083c6540022054d8d4206e206558e518d83c5740003c6640083c6840003c79400a205d18dc2066207d98ed58d82154d8d2330a17803c5b40383c5a40303c6c40383c6d40322054d8d4206e206558e518d83c5f40303c6e40383c6040403c71404a205d18dc2066207d98ed58d82154d8d2334a16603c5340383c5240303c6440383c6540322054d8d4206e206558e518d83c5740303c6640383c6840303c79403a205d18dc2066207d98ed58d82154d8d2330a16603c5b40283c5a40203c6c40283c6d40222054d8d4206e206558e518d83c5f40203c6e40283c6040303c71403a205d18dc2066207d98ed58d82154d8d233ca16403c5340283c5240203c6440283c6540222054d8d4206e206558e518d83c5740203c6640283c6840203c79402a205d18dc2066207d98ed58d82154d8d2338a16403c41400054931a8c9a403c4140093852400130501787d4697500000e780a080014903c524046306052003c5d40583c5c40503c6e40583c6f40522054d8d4206e206558e518d83c5140603c6040683c6240603c73406a205d18dc2066207d98ed58d82154d8d233ca14603c5540583c5440503c6640583c6740522054d8d4206e206558e518d83c5940503c6840583c6a40503c7b405a205d18dc2066207d98ed58d82154d8d2338a14603c5d40483c5c40403c6e40483c6f40422054d8d4206e206558e518d83c5140503c6040583c6240503c73405a205d18dc2066207d98ed58d82154d8d2334a14603c5540483c5440403c6640483c6740422054d8d4206e206558e518d83c5940403c6840483c6a40403c7b404a205d18dc2066207d98ed58d82154d8d2330a14603c5d40783c5c40703c6e40783c6f40722054d8d4206e206558e518d83c5140803c6040883c6240803c73408a205d18dc2066207d98ed58d82154d8d233ca13603c5540783c5440703c6640783c6740722054d8d4206e206558e518d83c5940703c6840783c6a40703c7b407a205d18dc2066207d98ed58d82154d8d2338a13603c5d40683c5c40603c6e40683c6f40622054d8d4206e206558e518d83c5140703c6040783c6240703c73407a205d18dc2066207d98ed58d82154d8d2334a13603c5540683c5440603c6640683c6740622054d8d4206e206558e518d83c5940603c6840683c6a40603c7b406a205d18dc2066207d98ed58d82154d8d2330a13683ca3404054b29a883ca340493854404130501467d4697400000e780205e014b03358179833501790336817883360178233ca15a2338b15a2334c15a2330d15a033501658335816503360166833681662338a126233cb1262330c1282334d128033501468335814603360147833681472334a1222338b122233cc1222330d124033581378335013703368136833601362338a1762334b1762330c176233cd1740335815b8335015b0336815a8336015a233ca1782338b1782334c1782330d178033501278335812703360128833681282338a164233cb1642330c1662334d166033581228335012303368123833601242338a172233cb1722330c1742334d174033501778335817603360176833681752330a172233cb1702338c1702334d170139a8903cee893f9790009456312a9041355ba03ac1a2e9503450500335535010589930a4008630a052c1305015a7d46814597400000e780803d88162c0b1306200497400000e7806049014a0149f1a1a28d230081469305017813060002130401781305114697400000e78020479305016513060002930401651305114897400000e780a045a300614b2301514b93050173130600021305314a97400000e780e04393058170130600021305314c97400000e780a0421355ba036e8aac1a2e95034505003355350105892c0b19e903498119034a91191304a1199304a11b9305114a03459401034684018346a4010347b4012205518dc2066207d98e558d0346d4018346c4010347e4018347f4012206558e4207e2075d8f598e0216518d233ca15a034514010346040183462401034734012205518dc2066207d98e558d034654018346440103476401834774012206558e4207e2075d8f598e0216518d2338a15a03459400034684008346a4000347b4002205518dc2066207d98e558d0346d4008346c4000347e4008347f4002206558e4207e2075d8f598e0216518d2334a15a034514000346040083462400034734002205518dc2066207d98e558d034654008346440003476400834774002206558e4207e2075d8f598e0216518d2330a15a03c5940003c6840083c6a40003c7b4002205518dc2066207d98e558d03c6d40083c6c40003c7e40083c7f4002206558e4207e2075d8f598e0216518d2330a17603c5140103c6040183c6240103c734012205518dc2066207d98e558d03c6540183c6440103c7640183c774012206558e4207e2075d8f598e0216518d2334a17603c5940103c6840183c6a40103c7b4012205518dc2066207d98e558d03c6d40183c6c40103c7e40183c7f4012206558e4207e2075d8f598e0216518d2338a17603c5140003c6040083c6240003c734002205518dc2066207d98e558d03c6540083c6440003c7640083c774002206558e4207e2075d8f598e0216518d233ca17488161306200497400000e780001f930a4008c669854d15a4034981199307a11903c5170083c5070003c6270083c6370022054d8d4206e206558e518d83c5570003c6470083c6670003c77700a205d18dc2066207d98ed58d82154d8d2330a15a03c5970083c5870003c6a70083c6b70022054d8d4206e206558e518d83c5d70003c6c70083c6e70003c7f700a205d18dc2066207d98ed58d82154d8d2334a15a03c5170183c5070103c6270183c6370122054d8d4206e206558e518d83c5570103c6470183c6670103c77701a205d18dc2066207d98ed58d82154d8d2338a15a03c5970183c5870103c6a70183c6b70122054d8d4206e206558e518d83c5d70103c6c70183c6e70103c7f701a205d18dc2066207d98ed58d82154d8d233ca15a9307a11b03c5970083c5870003c6a70083c6b70022054d8d4206e206558e518d83c5d70003c6c70083c6e70003c7f700a205d18dc2066207d98ed58d82154d8d2330a17603c5170183c5070103c6270183c6370122054d8d4206e206558e518d83c5570103c6470183c6670103c77701a205d18dc2066207d98ed58d82154d8d2334a17603c5970183c5870103c6a70183c6b70122054d8d4206e206558e518d83c5d70103c6c70183c6e70103c7f701a205d18dc2066207d98ed58d82154d8d2338a17603c5170083c5070003c6270083c6370022054d8d4206e20683c55700558e518d03c64700a20583c6670003c77700d18d034a9119c2066207d98ed58d82154d8d233ca174881613061002814597400000e78080efc66923042123a30441239305015a130600026a8597400000e780a0fa93058175130600025e8597400000e78080f9881c8c161306200497400000e78080f8630c0920281d0c041306100297400000e78040f703451d0083450d0003462d0083463d0022054d8d4206e206558e518d83455d0003464d0083466d0003477d00a205d18dc2066207d98ed58d82154d8d2330a17803459d0083458d000346ad008346bd0022054d8d4206e206558e518d8345dd000346cd008346ed000347fd00a205d18dc2066207d98ed58d82154d8d2334a17803451d0183450d0103462d0183463d0122054d8d4206e206558e518d83455d0103464d0183466d0103477d01a205d18dc2066207d98ed58d82154d8d2338a17803459d0183458d010346ad018346bd0122054d8d4206e206558e518d8345dd010346cd018346ed010347fd01a205d18dc2066207d98ed58d82154d8d233ca17803c59b0083c58b0003c6ab0083c6bb0022054d8d4206e206558e518d83c5db0003c6cb0083c6eb0003c7fb00a205d18dc2066207d98ed58d82154d8d233ca16403c51b0183c50b0103c62b0183c63b0122054d8d4206e206558e518d83c55b0103c64b0183c66b0103c77b01a205d18dc2066207d98ed58d82154d8d2330a16603c59b0183c58b0103c6ab0183c6bb0122054d8d4206e206558e518d83c5db0103c6cb0183c6eb0103c7fb01a205d18dc2066207d98ed58d82154d8d2334a16603c51b0083c50b0003c62b0083c63b0022054d8d4206e206558e518d83c55b0003c64b0083c66b0003c77b00a205d18dc2066207d98ed58d82154d8d2338a164054b95a01795feff9305c542130600021305912297400000e78000188345012701254d8d05e11795feff9305a540130600021305112797400000e780e01501256309055c281d0c041306100297400000e78000d2130501787d46ea8597400000e78000d1014be6e003450127630a05209307212703c5970183c5870103c6a70183c6b70122054d8d4206e206558e518d83c5d70103c6c70183c6e70103c7f701a205d18dc2066207d98ed58d82154d8d233ca14603c5170183c5070103c6270183c6370122054d8d4206e206558e518d83c5570103c6470183c6670103c77701a205d18dc2066207d98ed58d82154d8d2338a14603c5970083c5870003c6a70083c6b70022054d8d4206e206558e518d83c5d70003c6c70083c6e70003c7f700a205d18dc2066207d98ed58d82154d8d2334a14603c5170083c5070003c6270083c6370022054d8d4206e206558e518d83c5570003c6470083c6670003c77700a205d18dc2066207d98ed58d82154d8d2330a1469307212903c5970083c5870003c6a70083c6b70022054d8d4206e206558e518d83c5d70003c6c70083c6e70003c7f700a205d18dc2066207d98ed58d82154d8d2334a13603c5170183c5070103c6270183c6370122054d8d4206e206558e518d83c5570103c6470183c6670103c77701a205d18dc2066207d98ed58d82154d8d2338a13603c5970183c5870103c6a70183c6b70122054d8d4206e206558e518d83c5d70103c6c70183c6e70103c7f701a205d18dc2066207d98ed58d82154d8d233ca13603c5170083c5070003c6270083c6370022054d8d4206e206558e518d83c5570003c6470083c6670003c77700a205d18dc2066207d98ed58d8215034911274d8d2330a136854c29a803491127130501467d469305212797400000e780e0ad814c03358179833501790336817883360178233ca1342338b1342334c1342330d134033501658335816503360166833681662330a1322334b1322338c132233cd132033501468335814603360147833681472330a1302334b1302338c130233cd13003358137833501370336813683360136233ca12e2338b12e2334c12e2330d12e63030c028a642c1d62859770ffffe780c0ba2e8471c5638604120e046294033c8472fd14cdb7900508622330a15608660c6a030686018334812b2334a1562338b156230cc1569770ffffe780809f833501562a84233c955a033581562330b45c83350157233004002334a45c030581572338b45c8544231b945a230ca45c23046401a30444011305a4008c061306000297400000e780409c1305a4020c161306000297400000e780209b23059405a30524051305c4040c061306000297400000e78080991305c4068c151306000297400000e7806098a2fc02e1866c6f001002330554032a9c23046c01a3044c011305ac008c061306000297400000e780c0951305ac020c161306000297400000e780a09423059c05a3052c051305cc040c061306000297400000e78000931305cc068c151306000297400000e780e091866c7daf4afc940588628c66906a83c686012330a1562334b1562338c156230cd156230cd1582338c1582334b1582330a15883596c5b0339812b2d4563f9a906da8dd28b13058c5b130b140093145400b3058500ae94330a540363fc69072380240113558903a383a400135509032383a40013558902a382a400135509022382a40013558901a381a400135509012381a40013558900a380a4001385840093050158654697400000e78020876da0930b4008054d914a154552f85af46369a4126303a412014d19456311a4120144954a39aa93155b005a952e9533848940131654002296a68597400000e780e0c713558903a383a400135509032383a40013558902a382a400135509022382a40013558901a381a400135509012381a40013558900a380a400238024011385840093050158654697300000e780207e13058c00b305450133065b0332953306540397400000e78060c18529629a2304ba01a3047a011305aa008c061306000297300000e780a07a1305aa020c161306000297300000e780807923059a056275a305aa041305ca040c061306000297300000e780c0771305ca068c151306000297300000e780a076231b3c5b854d6da463020c600a653384ad400c0462859770ffffe780e08a630f05586305b45f8e05e29503bc85720504cdb7a28a19a06514994a9760ffffe78020712a8b23300500231b055a83596c5b93c4faffce94231b955a930d8c5b93955a0033855d01aa95130501651306100297300000e780206f130a8c0033857a035295834b050093051500130501781306300897300000e780006d314563e4a4006f10a06c66f0ea8c138d1a003385a941630495006f10e07213058b5b93155d00ea9dee9513965400269697300000e780806913064008b305cd02d29513058b003386c40297300000e780e067231b5c5b1305015a930501651306100297300000e780606613050146930501781306300897300000e7802065628d63930c005a8d83596d5b13058d5b930d140093145400b3058500ae94930a4008330a540363fab9052380240113558903a383a400135509032383a40013558902a382a400135509022382a40013558901a381a400135509012381a40013558900a380a4001385840093050158654697300000e780a05d59a093955d006e952e9533848940131654002296a68597400000e780a0a013558903a383a400135509032383a40013558902a382a400135509022382a40013558901a381a400135509012381a40013558900a380a400238024011385840093050158654697300000e780e05613058d00b305450133865d0332953306540397400000e780209a854d027485296a9a22752304aa004275a304aa001305aa008c061306000297300000e780e0521305aa020c161306000297300000e780c05123058a046275a305aa041305ca040c061306000297300000e78000501305ca068c151306000297300000e780e04e231b3d5b130581759305015a1306100297300000e780604d8816930501461306600897300000e780404c130da12209456397ab00930ba124866cc669b9a613058162930581751306100297300000e780c0491305015a8c161306300897300000e780a04803350c00c669014a630705225a84835c4c5b2a8c13058170930581621306100297300000e7802046230071479305015a130630081305114697300000e780a044630400006f10804783596c5b2d4563eba92a52fc854d114a154522f8930b400863efac006389ac00814d19456397ac00814c154a29a0668a19a0e51c194a9760ffffe78060412a8b23300500231b055a03596c5b9344faffca94231b955a930a8c5b93155a0033854a01aa95130581751306100297300000e780e03c13048c0033057a032295034d05009305150088161306300897300000e780e03a314563e4a4006f10803aee8b930d1a003305b941630495006f10603d13058b5b93955d00ee9ad69513965400269697300000e7808037930a4008b3855d03a29513058b003386540397300000e780e035231b4c5b13050173930581751306100297300000e7806034130501788c161306300897300000e780403303546b5b13051400b1456364b4006f10c032338649416304a6006f104036627a050a8e0de29d93858d7293048b720e06268597300000e780a02f014593153500a6958c6133368500239aa55a3295b336a40093c61600758e23b0650165f21305016e930501731306100297300000e780202c13050165930501781306300897300000e780e02a6285854dc66963930b005a851306817093060146e68542779760ffffe780802c0945630fad10ea8b130581629305016e1306100297300000e78020271305015a930501651306300897300000e780e02503350c005a84e31e05dce67499e06f10e02d0a699760ffffe78040252a8423300500231b055a233495721305190080e0239a045aa2fc2ae1130da122866c630449016f10402b8354645b2945637495006f10402b130984721b851400231ba45a13955400b30594002e951305855b930581621306100297300000e780001e3385540322952304750125059305015a1306300897300000e780401c8504139534004a952330650123308b00231a9b5aa1a02300015a631eb40923308137233401362338b136130501468c161306015a9760ffffe780203559aa13068170930601466285e68522879760ffffe780a01ac669130da122866c930ba124aa64850426e57e75de753e769e762aeb2ee732e3b6fe280b90133414981cce8597a0ffffe780009d13f51c00631e0516a66413f5f40f130515f0933c1500138414008813ac1a26869750ffffe780c0e3a6896fe0afe18e05e29503b5857219c8b30580400356655b0e06329503358572fd15edf98355655bfd152338a164233c01642330b16613050146930501651306015a9760ffffe780402913050178930501461306500a97300000e780600b03358150033a81518355655b03340151aa84636fba00046191c8035a455b83d5645b05042685e378bafe19a0228a2a8413155a00b38544012e959309855b33055a03269513098500881613061002ce8597300000e780e00593050178130610024e8597300000e780c0041306400813051138ca8597300000e780a003130640084a859305117a97300000e780800209cc0e0ad29483b404737d14c66919c483b484727d146dfc11a0c669130501468c161306500a97300000e780a0ff23349150233801502a658345015a7d152ae5e38505e8667519e16f10200c8a6599e16f10400c03368572b2fcfd152ee12330060097f0feffe78000ad85b5a8082c0b97a0ffffe78000a16fd00ff92689aa84033a8148833a014813155900229583459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18d233cb13683451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2338b13683459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2334b13683451500034605008346250003473500a205d18dc20662070346550083474500d98ed58d22065d8e834665000347750093174900b309f400c2066207d98e558e0216d18d2330b136930501781306000297300000e78020e803b5891683b5091623b0591723b4491791cc0e094a9403348422fd14930a400881c803340422fd14edfc19a0930a400803368137833601370337813683370136233cc1462338d1462334e1462330f1462330b1482334a14823388148233c01480a758345015a7d152af199e16fe0afad4a65e30d0570ea65e38f05700336052232e9fd152eed2338062097f0feffe78020906fe04fabe6650676a6762eef467732f336f7e6753afb2a660a643339b000b3062041b3f9c600638d09063336200193361500758e11ca054909c483b585727d146dfc014a2e8521a02e8ae30a09668355655b6362b4020461e381045a0354455b050a97f0feffe780808983d5645b2685e373b4fe26858145fd190504e3050afa0e042295033585729304faff81450144d9d803358572fd14edfc8145014461b7630a090219e52e8509c4033585727d146dfc0c6191c92e8497f0feffe78020840c602285edf911a02a84228597f0feffe780e082ca6501450a766a6a3339b000b3062041b3f9c600638e09063336200193361500758e01ce054963070a0083b505227d1ae31d0afe81442e8521a0ae84e30c095a8355a5216363ba0203340521e306044e035a8521850497e0feffe780007d8355a4212285e372bafe22858145fd19050ad5d00e0a529503350522fd148145014ad1d803350522fd14edfc8145014a59b7630e090209e92e8563070a00033505227d1ae31d0afe8335052199c92e8497e0feffe7808077833504212285e5f911a02a84228597e0feffe780207613050004854597e0feffe780c074e3040558aa8dc26703c5970183c5870103c6a70183c6b70122054d8d4206e206558e518d83c5d70103c6c70183c6e70103c7f701a205d18dc2066207d98ed58d82154d8d233ca14603c5170183c5070103c6270183c6370122054d8d4206e206558e518d83c5570103c6470183c6670103c77701a205d18dc2066207d98ed58d82154d8d2338a14603c5970083c5870003c6a70083c6b70022054d8d4206e206558e518d83c5d70003c6c70083c6e70003c7f700a205d18dc2066207d98ed58d82154d8d2334a14603c5170083c5070003c6270083c6370022054d8d4206e206558e518d83c5570003c6470083c6670003c77700a205d18dc2066207d98ed58d82154d8d2330a146130501482c0b1306000297300000e78080b293050146130600046e8597300000e78060b185458546854c6e8501469770ffffe780409d6265033c050109452afa02fe82e2e3090c280949014b014482e46265033a05001785feff1305e598aae893044006130d00108949b3058a0003c50500130685fba546e3eec62a0e06c66636961062930a14000286e36f2b23d27933059b024e950344e5fb130940068944e307943e1306c5f9835bc5f90355c6018355a6018356e6010357060242054d8d82164217d98e558d2334a1280355460183552601835666010357860142054d8d82164217d98e558d2330a1280355c6008355a60042058356e600035706014d8d9305360282164217d98e558d233ca126035546008356260003576600035686004205558d02174216598e518d2338a126130610041305117897300000e780a09f23008178791bdae233052b034e95034425020949e3029434835405008355c5010356a5018356e50103570502c205d18d82164217d98ed58daee183554501035625018356650103578501c205d18d82164217d98ed58d2efd8355c5000356a500c2058356e500035705014d8e9305350282164217d98e558e32f9035645008356250003576500035585004206558e02174215598d518d2af5130610041305113697300000e780209533c574011335150093b50b106d8d23008136e307050ca8082c115e869740ffffe78060651305015a8c1c5e869740ffffe7806064a8089305015a1306000297300000e78040d30125e31c050813958b036d912c112e950345050093f57b003355b5000589630d056c13050146b008930601789816d9ad2665e314050626651a056e9583459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18d233cb14683451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2338b14683459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2334b14683451500034605008346250003473500a205d18dc2066207d98ed58d034655008346450003476500834775002206558e4207e2075d8f598e0216d18d2330b14683459503034685038346a5030347b503a205d18dc2066207d98ed58d0346d5038346c5030347e5038347f5032206558e4207e2075d8f598e0216d18d233cb13683451503034605038346250303473503a205d18dc2066207d98ed58d034655038346450303476503834775032206558e4207e2075d8f598e0216d18d2338b13683459502034685028346a5020347b502a205d18dc2066207d98ed58d0346d5028346c5020347e5028347f5022206558e4207e2075d8f598e0216d18d2334b13683451502034605028346250203473502a205d18dc2066207d98ed58d034655028346450203476502034575022206558e42076205598df276518d02154d8d2330a1366319db00081ada859790ffffe78040ec166bd27933059b023384a9002310040013052400930501461306000297200000e780a06923010402130534028c161306000297200000e7804068050bdae226650505aae4f9a133356001b3b58a016d8d630e055ed29a83ca0a0063940a00930a00107d1bdae233059b024e9583442502638b247b835c05008355c5010356a5018356e50103570502c205d18d82164217d98ed58d233cb13683554501035625018356650103578501c205d18d82164217d98ed58d2338b1368355c5000356a500c2058356e500035705014d8e9305350282164217d98e558e2334c136035645008356250003576500035585004206558e02174215598d518d2330a136130501461306100497200000e780205b03358137833501370336813683360136aaf8aef4b2f0b6ec2300917893050146130610041305117897200000e780205863f7ac514675a6750676e666233ca15a2338b15a2334c15a2330d15a63820a2c8144b38b9c0013950b0341916371a54f1305015aac085e869740ffffe780a02613958b036d91ac082e950345050093f57b003355b500058915c11305014613061002814597200000e780804488161306015a93060146130701780da01305014613061002814597200000e780604288161306015a9306017813070146de859790ffffe78000d78504130501788c161306200497200000e780804c139504034191e36155f739ac63050b44930b140263e48b50636f7c43637f746133855b4193050002631eb55cb3055a01130600021305117897200000e78080487d1bdae2d2792300017833059b024e958344250289456392b408dda3630d0b3e930b240463e18b4c63677c3f63f38a4d130524026360ac4c63e2ab5c130940063386ab4093060002631ed656d29a83c40a0013842500b305aa00130600021305217a97200000e780e0411306000213052178a28597200000e780c0407d1bdae2d279a30091782300917933052b034e95834425028945638ab456035405008355c5010356a5018356e50103570502c205d18d82164217d98ed58daef883554501035625018356650103578501c205d18d82164217d98ed58daef48355c5000356a500c2058356e500035705014d8e9305350282164217d98e558eb2f0035645008356250003576500035585004206558e02174215598d518daaec130610041305113697200000e780e035230091366374a42f1305015aac0822869740ffffe780e006131584036d91ac082e9503450500937574003355b500058909c9130501461306015a93060178981601a8130501461306015a941613070178a2859790ffffe78080b9930440067275631cab000949081ada859790ffffe78020af166bd27911a00949050433059b02b384a90023908400138524009305015a1306000297200000e780202c1385240293044006930501461306200497200000e780a02a050bdae2de8ae5a8e68b0335015a8335815a0336015b8336815b2330a1362334b1362338c136233cd13613050146930501781306200497200000e780c0267275631aab00081ada859790ffffe78000a6166bd279854c93044006930a2400850b33059b023384a90023107401130524008c161306000297200000e780c02213052402930501461306200497200000e7808021166b9da013050146b008941613070178de859790ffffe78020a9930440067275631aab00081ada859790ffffe780e09e166bd279850b33059b023384a9002310740113052400ac081306000297200000e780401c13052402930501461306200497200000e780001b050bdae2568463ed8aed05456319ab1252740355040013450510a66593c515004d8d631e051093052402130511659790ffffe780a0bd727511c5228597e0feffe780e0c76e8597e0feffe78040c703156165831541650356216583061165231aa172c205d18d033581662328b1728305016703348165233ca174833401662300b1762304d1221305912293050173194697200000e780801113558403230ba12213550403a30aa12213558402230aa12213550402a309a122135584012309a12213550401a308a122135584002308a122a307812213d58403230fa12213d50403a30ea12213d58402230ea12213d50402a30da12213d58401230da12213d50401a30ca12213d58400230ca122a30b91221305f12393058175254697200000e780e008281413060002a26597200000e780604a814c01251334150005a0854c727511c5527597e0feffe78060b76e8597e0feffe780c0b613044002e265886511c5886197e0feffe78080b56685a2850d618330817e0334017e8334817d0339017d8339817c033a017c833a817b033b017b833b817a033c017a833c8179033d0179833d81781301017f8280a308a16441bfad452685ada0b1459da097e0feffe78000b01775feff1305a56c09a897e0feffe780e0ae1775feff1305856b9305b00291a81785feff130515839305500399a01775feff1305b57f25a81775feff1305157f3da01775feff1305656b29a01775feff1305c56af14531a85685e2859730ffffe78040f500001775feff1305357c930580029720ffffe780a06900001775feff1305e56459bf1775feff1305257593050003c5b71775feff1305655f93050002c9bfad4566855dbf1775feff130515787dbf1775feff1305757755bf1775feff1305e56099bf1775feff13054560b1b71775feff1305a55f89b71775feff1305e5729305100271b7ad454e8585bf1775feff1305b573a5bf1775feff1305255d29bf1775feff13056570e1bf1775feff1305e55b19b71775feff1305256c85bf1775feff1305a55695bf13050002930500022db71305000497e0feffe780809d00001775feff13058558c1bd1775feff1305e557d9b51775feff1305455775bd5685de85e5bd1775feff1305455675b51775feff1305a5554db5034715008347050022075d8f83472500c207d98f0347350062075d8f834745008217d98f0347550022175d8f8347650003457500c217d98f62155d8d82802e869737000083b7675c814582870971a2faa6f6caf286feceeed2ead6e6dae25efe62fa66f66af26eee2ae4ae8401441309000833858400eff0bff8930704018a9788e32104e31724ffa265130600040809ef10d05d4a754a6fc2679782feff83b242942a9f3e9fa267e269ea78b4639787feff83b78795ea6eb346df00bd8e939706028192dd8eb692334555009357850122155d8d4e9f2a9fb346df0093d70601c216dd8eb69233c5a200931715007d915d8d8277c69e978ffeff83bf0f90be9ea2670e660a7eb8679787feff83b7678ec27b33c7ee003d8f9317070201935d8fba9fb3c8f80193d78801a218b3e8f800a277329e5e9ebe9ec69e33c7ee009357070142175d8fba9fb3c81f019397180093d8f803b3e8f800a2679785feff83b5c58b978cfeff83bc4c88bc6b2e682a73b347fe00ad8f939507028193cd8fbe9c334696019355860122164d8ee275066442932e9e329eb347fe0093d50701c217cd8fbe9c33c6cc00931516007d924d8ea26522939783feff83b3a384ac6d178dfeff033d0d85a664b345b300b3c57500939305028191b3e575002e9d3348a80193538801221833687800269342934669b345b30093d30501c215b3e575002e9d4a9f33480d01469f93131800b345bf001358f80333687800939305028191b3e57500666bae9cb3c81c0193d38801a218b3e878005a9f469f067ab345bf0093d30501c215b3e57500ae9cd29eb3c81c01b29e93931800b3c6de0093d8f803b3e87800939306028192b3e67600a674369d3346cd0093538601221633667600a69eb29eb3c6de0093d30601c216b3e67600369d3346cd00931316007d9233667600c673e67a0a6c1e9e429e3347ee00931407020193458fba9233c8020193548801221833689800569e429e3347ee00935407014217458fba92629333c802012a9393141800b347f3001358f80333689800939407028193c58fbe9f33c5af00935485012215458daa64629fde9e26932a93b347f30093dd0701c217b3e7b701be9f33c5af00931d15007d913365b5012a9fb346df00939d06028192b3e6b601b69233c5a200935d850122153365b501529f2a9fb346df0093dd0601c216b3e6b601b69233c5a200c69e931d150033c7ee007d913365b501931d070201933367b701ba9fb3c81f0193dd8801a218b3e8b801ca9ec69e33c7ee00935d070142173367b701ba9f5a9eb3c81f01329e939d1800b347fe0093d8f803b3e8b801939d07028193b3e7b701be9c33c6cc00935d860122163366b601269e329eb347fe0093dd0701c217b3e7b701be9c569333c6cc004293931d1600b345b3007d923366b601939d05028191b3e5b5012e9d33480d01935d880122183368b80122934293b345b30093dd0501c215b3e5b5012e9d4e9f33480d01469f931d1800b345bf001358f8033368b801939d05028191b3e5b501ae9cb3c81c0193dd8801a218b3e8b8011e9f469fb345bf0093dd0501c215b3e5b501ae9cb3c81c01939d180093d8f803b3e8b801c26dee9eb29eb3c6de00939d06028192b3e6b601369d3346cd00935d860122163366b601827dee9eb29eb3c6de0093dd0601c216b3e6b601369d3346cd00931d16007d923366b601a67d9e9ec69e6e9e429e3347ee00931d070201933367b701ba9233c80201935d880122183368b801a66d6e9e429e3347ee00935d070142173367b701ba9233c80201931d18001358f8033368b801e27d33c7ee006e932a93b347f300939d07028193b3e7b701be9f33c5af00935d850122153365b501a27d6e932a93b347f30093dd0701c217b3e7b701be9f33c5af00931d15007d913365b501a67d269342936e9f2a9fb346df00939d06028192b3e6b601b69233c5a200935d850122153365b5014a9f2a9fb346df0093dd0601c216b3e6b601b69233c5a200931d15007d913365b501931d070201933367b701ba9fb3c81f0193dd8801a218b3e8b801c26db345b3005693ee9ec69e33c7ee00935d070142173367b701ba9fb3c81f01939d180093d8f803b3e8b801e27d529f469f6e9e329eb347fe00939d07028193b3e7b701be9c33c6cc00935d860122163366b601827d6e9e329eb347fe0093dd0701c217b3e7b701be9c33c6cc00931d16007d923366b601939d05028191b3e5b5012e9d33480d01935d880122183368b8014293b345b30093dd0501c215b3e5b5012e9d33480d01931d1800b345bf001358f8033368b801939d05028191b3e5b501ae9cb3c81c0193dd8801a218b3e8b801629f469fb345bf0093dd0501c215b3e5b501ae9cb3c81c01939d180093d8f803b3e8b801a27d5a932a93ee9eb29eb3c6de00939d06028192b3e6b601369d3346cd00935d860122163366b601a29eb29eb3c6de0093dd0601c216b3e6b601369d3346cd00931d16007d923366b601a66db347f3005e936e9e429e3347ee00931d070201933367b701ba9233c80201935d880122183368b8014e9e429e3347ee00935d070142173367b701ba9233c80201931d18001358f8033368b801939d07028193b3e7b701be9f33c5af00935d850122153365b5012a93b347f30093dd0701c217b3e7b701be9f33c5af00931d15007d913365b501a66d569e329e6e9f2a9fb346df00939d06028192b3e6b601b69233c5a200935d850122153365b5015a9f2a9fb346df0093dd0601c216b3e6b601b69233c5a200931d15007d913365b501a27db347fe001e9eee9ec69e33c7ee00931d070201933367b701ba9fb3c81f0193dd8801a218b3e8b801ce9ec69e33c7ee00935d070142173367b701ba9fb3c81f01939d180093d8f803b3e8b801939d07028193b3e7b701be9c33c6cc00935d860122163366b601329eb347fe0093dd0701c217b3e7b701be9c33c6cc00931d16007d923366b601a67d5e9e6e934293b345b300939d05028191b3e5b5012e9d33480d01935d880122183368b80162934293b345b30093dd0501c215b3e5b5012e9d33480d01931d18001358f8033368b801827d429e3347ee006e9f469fb345bf00939d05028191b3e5b501ae9cb3c81c0193dd8801a218b3e8b801229f469fb345bf0093dd0501c215b3e5b501ae9cb3c81c01939d180093d8f803b3e8b801e27d26932a93ee9eb29eb3c6de00939d06028192b3e6b601369d3346cd00935d860122163366b601d29eb29eb3c6de0093dd0601c216b3e6b601369d3346cd00931d16007d923366b601931d070201933367b701ba9233c80201935d880122183368b801c26db347f3004a936e9e429e3347ee00935d070142173367b701ba9233c80201931d18001358f8033368b801939d07028193b3e7b701be9f33c5af00935d850122153365b5012a93b347f30093dd0701c217b3e7b701be9f33c5af00931d15007d913365b5015a9f2a9fb346df00939d06028192b3e6b601b69233c5a200935d850122153365b501c26d529342936e9f2a9fb346df0093dd0601c216b3e6b601b69233c5a200931d15007d913365b501e27db345b3002693ee9ec69e33c7ee00931d070201933367b701ba9fb3c81f0193dd8801a218b3e8b801a66d629fee9ec69e33c7ee00935d070142173367b701ba9fb3c81f01939d180093d8f803b3e8b801827d469f6e9e329eb347fe00939d07028193b3e7b701be9c33c6cc00935d860122163366b6015e9e329eb347fe0093dd0701c217b3e7b701be9c33c6cc00931d16007d923366b601939d05028191b3e5b5012e9d33480d01935d880122183368b8014293b345b30093dd0501c215b3e5b5012e9d33480d01931d1800b345bf001358f8033368b801939d05028191b3e5b501ae9cb3c81c0193dd8801a218b3e8b8014e9f469fb345bf0093dd0501c215b3e5b501ae9cb3c81c01939d180093d8f803b3e8b801a67d229e429eee9eb29eb3c6de00939d06028192b3e6b601369d3346cd00935d860122163366b6019e9eb29eb3c6de0093dd0601c216b3e6b601369d3346cd00931d16003347ee007d923366b601931d070201933367b701ba9233c80201935d880122183368b8014a9e429e3347ee00935d070142173367b701ba9233c80201931d18001358f8033368b801a27da29ec69e6e932a93b347f300939d07028193b3e7b701be9f33c5af00935d850122153365b50156932a93b347f30093dd0701c217b3e7b701be9f33c5af00931d15007d913365b501827d33c7ee00d29e6e9f2a9fb346df00939d06028192b3e6b601b69233c5a200935d850122153365b5011e9f2a9fb346df0093dd0601c216b3e6b601b69233c5a200931d15007d913365b501931d070201933367b701ba9fb3c81f0193dd8801a218b3e8b801c69e33c7ee00935d070142173367b701ba9fb3c81f01939d180093d8f803b3e8b801c26d4a9342936e9e329eb347fe00939d07028193b3e7b701be9c33c6cc00935d860122163366b601a67db345b3005e9f6e9e329eb347fe0093dd0701c217b3e7b701be9c33c6cc00931d16007d923366b601939d05028191b3e5b5012e9d33480d01935d880122183368b801a27d469f269e6e934293b345b30093dd0501c215b3e5b5012e9d33480d01931d1800b345bf001358f8033368b801939d05028191b3e5b501ae9cb3c81c0193dd8801a218b3e8b801569f469fb345bf0093dd0501c215b3e5b501ae9cb3c81c01939d180093d8f803b3e8b801a66d429e3347ee00ee9eb29eb3c6de00939d06028192b3e6b601369d3346cd00935d860122163366b601e27d629e4e93ee9eb29eb3c6de0093dd0601c216b3e6b601369d3346cd00931d16007d923366b601931d070201933367b701ba9233c80201935d880122183368b801429e3347ee00935d070142173367b701ba9233c802012a93931d1800b347f3001358f8033368b801939d07028193b3e7b701be9f33c5af00935d850122153365b5015a932a93b347f30093dd0701c217b3e7b701be9f33c5af00931d15007d913365b5011e9f2a9fb346df00939d06028192b3e6b601b69233c5a200935d850122153365b501e27dce9ec69e6e9f2a9fb346df0093dd0601c216b3e6b601b69233c5a200931d150033c7ee007d913365b501931d070201933367b701ba9fb3c81f0193dd8801a218b3e8b801a69ec69e33c7ee00935d070142173367b701ba9f629eb3c81f01329e939d1800b347fe0093d8f803b3e8b801939d07028193b3e7b701be9c33c6cc00935d860122163366b601569e329eb347fe0093dd0701c217b3e7b701be9c5e9333c6cc004293931d1600b345b3007d923366b601939d05028191b3e5b5012e9d33480d01935d880122183368b80152934293b345b30093dd0501c215b3e5b5012e9d33480d01931d18001358f8033368b801c26da29eb29e6e9f469fb345bf00939d05028191b3e5b501ae9cb3c81c0193dd8801a218b3e8b801a66db3c6de005a9e6e9f469fb345bf0093dd0501c215b3e5b501ae9cb3c81c01939d180093d8f803b3e8b801939d06028192b3e6b601369d3346cd00935d860122163366b601a27d429e3347ee00ee9eb29eb3c6de0093dd0601c216b3e6b601369d3346cd00931d16007d923366b601931d070201933367b701ba9233c80201935d880122183368b801827d4a932a936e9e429e3347ee00935d070142173367b701ba9233c80201931d1800b347f3001358f8033368b801939d07028193b3e7b701be9f33c5af00935d850122153365b501a67d569f1e9e6e932a93b347f30093dd0701c217b3e7b701be9f33c5af00931d15007d913365b5012a9fb34ddf0093960d0293dd0d02b3eddd00ee92b3c6a20013d58601a216c98e2675329eb347fe002a9f369fb34dbf0113d50d01c21db3edad00ee92b3c6d20013951600fd92c98e26654e9eaa9ec69e33c7ee00131507020193498fba9fb3c81f0113d58801a218b3e8a800e29ec69e33c7ee00135507014217498fba9fb3c81f011395180093d8f803b3e8a800139507028193c98fbe9c33c6cc00135586012216498e329eb347fe0013d50701c217c98fbe9c33c6cc00131516007d92498e2275a69eb29e2a934293b345b300139505028191c98d2e9d33480d011355880122183368a8005a934293b345b30013d50501c215c98d2e9d33480d01131518001358f8033368a8006275b3cdbe01de9e2a9f469fb345bf00139505028191c98dae9cb3c81c0113d58801a218b3e8a80042654a9e429e2a9f469fb345bf0013d50501c215c98dae9cb3c81c011395180093d8f803b3e8a80013950d0293dd0d02b3edad006e9d3346cd00135586012216498eb29eb3cdbe0113d50d01c21db3edad006e9d3346cd00131516003347ee007d92498e131507020193498fba9233c802011355880122183368a800229e429e3347ee00135507014217498fba9233c80201131518001358f8033368a8000275229fe29e2a933693b347f300139507028193c98fbe9fb3c6df0013d58601a216c98e52933693b347f30013d50701c217c98fbe9fb3c6df0013951600fd92c98e369fb34dbf0113950d0293dd0d02b3edad00ee92b3c6d20013d58601a216c98e269f369fb34dbf0113d50d01c21db3edad00ee92b3c6d200c69e1395160033c7ee00fd92c98e131507020193498fba9fb3c81f0113d58801a218b3e8a800da9ec69e33c7ee00135507014217498fba9fb3c81f011395180093d8f803b3e8a80026751e9f469f2a9e329eb347fe00139507028193c98fbe9c33c6cc00135586012216498e2275d69e2a9e329eb347fe0013d50701c217c98fbe9c33c6cc00131516007d92498e4265b29eb3cdbe012a934293b345b300139505028191c98d2e9d33480d011355880122183368a8004a934293b345b30013d50501c215c98d2e9d33480d0113151800b345bf001358f8033368a800139505028191c98dae9cb3c81c0113d58801a218b3e8a80002754e9e429e2a9f469fb345bf0013d50501c215c98dae9cb3c81c011395180093d8f803b3e8a80013950d0293dd0d02b3edad006e9d3346cd00135586012216498e26653347ee005e9eaa9eb29eb3cdbe0113d50d01c21db3edad006e9d3346cd00131516007d92498e131507020193498fba9233c802011355880122183368a800429e3347ee00135507014217498fba92529333c80201369313151800b347f3001358f8033368a800139507028193c98fbe9fb3c6df0013d58601a216c98e6275529fca9e2a933693b347f30013d50701c217c98fbe9fb3c6df0013951600fd92c98e369fb34dbf0113950d0293dd0d02b3edad00ee92b3c6d20013d58601a216c98e0275c69e33c7ee002a9f369fb34dbf0113d50d01c21db3edad00ee92b3c6d20013951600fd92c98e131507020193498fba9fb3c81f0113d58801a218b3e8a800de9ec69e33c7ee00135507014217498fba9fb3c81f011395180093d8f803b3e8a80026654e9342932a9e329eb347fe00139507028193c98fbe9c33c6cc00135586012216498e229e329eb347fe0013d50701c217c98fbe9c33c6cc0013151600b345b3007d92498e139505028191c98d2e9d33480d011355880122183368a8006275269f469f2a934293b345b30013d50501c215c98d2e9d33480d0113151800b345bf001358f8033368a800139505028191c98dae9cb3c81c0113d58801a218b3e8a8002675da9eb29e2a9f469fb345bf0013d50501c215c98dae9cb3c81c0113951800b3cdbe0193d8f803b3e8a80013950d0293dd0d02b3edad006e9d3346cd00135586012216498ee29eb29eb3cdbe0113d50d01c21db3edad006e9d3346cd00131516007d92498e2275569336932a9e429e3347ee00131507020193498fba9233c802011355880122183368a8001e9e429e3347ee00135507014217498fba9233c8020113151800b347f3001358f8033368a800139507028193c98fbe9fb3c6df0013d58601a216c98e42655e9e329e2a933693b347f30013d50701c217c98fbe9fb3c6df0013951600fd92c98e4265b347fe0022932a9f369fb34dbf0113950d0293dd0d02b3edad00ee92b3c6d20013d58601a216c98e4e9f369fb34dbf0113d50d01c21db3edad00ee92b3c6d20013951600fd92c98e02754293b345b300aa9ec69e33c7ee00131507020193498fba9fb3c81f0113d58801a218b3e8a80022754a9faa9ec69e33c7ee00135507014217498fba9fb3c81f011395180093d8f803b3e8a800139507028193c98fbe9c33c6cc00135586012216498e6275469fd29e2a9e329eb347fe0013d50701c217c98fbe9c33c6cc00131516007d92498e139505028191c98d2e9d33480d011355880122183368a8002665b29eb3cdbe012a934293b345b30013d50501c215c98d2e9d33480d0113151800b345bf001358f8033368a800139505028191c98dae9cb3c81c0113d58801a218b3e8a8005a9f469fb345bf0013d50501c215c98dae9cb3c81c011395180093d8f803b3e8a80013950d0293dd0d02b3edad006e9d3346cd00135586012216498e26751e9e429eaa9eb29eb3cdbe0113d50d01c21db3edad006e9d3346cd00131516003347ee007d92498e131507020193498fba9233c802011355880122183368a800569e429e3347ee00135507014217498fba92629333c80201369313151800b347f3001358f8033368a800139507028193c98fbe9fb3c6df0013d58601a216c98e26933693b347f30013d50701c217c98fbe9fb3c6df0013951600fd92c98e7a9c369cb34dbc0113950d0293dd0d02b3edad00ee92b3c6d20013d58601a216c98e629a369ab34dba0113d50d01c21db3edad00ee92f69bb3c6d200c69b1395160033c7eb00fd92c98e131507020193498fba9fb3c81f0113d58801a218b3e8a8005e9946993347e900135507014217498fba9f729bb3c81f01329b13951800b347fb0093d8f803b3e8a800139507028193c98fbe9c33c6cc00135586012216498eda94b294a58f13d50701c217c98fbe9c9a9a33c6cc00c29a13151600b3c5ba007d92498e139505028191c98d2e9d33480d011355880122183368a80056944294a18d13d50501c215c98d2e9dd29933480d01c69913151800b3c5b9001358f8033368a800139505028191c98dae9cb3c81c0113d58801a218b3e8a800ce93c6931ee9b3c3b30093d50301c213b3e3b3009e9ce6f1b3cc1c0193951c0093dcfc03b3e595012efdc2651ee6ca95b295b3cdb50113950d0293dd0d02b3edad006e9d3346cd00135586012216498e0275aa95b2952eedb3c5b50113d50501c215c98d2e9deaf5334dcd0013161d00135dfd033366a601b2e12676aef926964296318f1315070293550702c98dae9233c802011357880122183368e8002667329742973af12d8f135607014217518fba9296e9b3c20201bafd1397120093d2f20333675700bae5627722973697b98f9395070213d607024d8eb29fb3c6df0093d78601a216dd8ea277ba97b6973ef5b18f13d70701c217d98fbe9ffeedb3cfdf003ee293971f0093dfff03b3e7f7013ef9a26714091386070498638c62a107a1062d8f8c7e2d8f23bce7fee317f6fef6705674b6741679f669566ab66a166bf27b527cb27c127df26d19618280397156e4833a050e52e8130a000822f826f44af04eec06fc330a5a412a842e89b284930905066373ca0452862330050e33855901ef00a0323c603864938404f8938707083ce093b70708ba9752993ce4ce852285d694efe08fceb30a9900130a0008b3859a402e8963649a0268702686ca854e95ef00a02e7c70e2700279a6977cf04274a274e269426aa26a216182803c6038642285938707083ce093b70708ba973ce4efe0afc9938404f85dbf797122f04ae82a842e891306800b81451305050426ec4ee406f4ef00801c9767feff83b747e01ce09767feff83b727e11ce49767feff83b787df1ce89767feff83b767e11cec9767feff83b747e01cf09767feff83b727de1cf49767feff83b707e01cf89767feff83b7e7dd1cfc81449309000433059900efe0cfbc330794001c63a104a98f1ce3e39634ff83470900a270e2647cf402744269a269014545618280357122e926e54ae106ed2a84b2843689eff0fff4634805021306000881450a85ef0000124a86a6850a85ef00401e8a85228513060008eff0bfe7930500080a85efe00fbaea604a64aa640a6901450d61828009ca411106e4eff09fe5a260014541018280014582801d71a2e8a6e4cae02a84ae843289814513068003280086ec02e0ef00e00b7d55d5c47c747d556363f90a3c68c5e368703c603864aa973ce0b3b7a700ba973ce48347040f99c3fd573cecfd571309040613060008098e3ce881454a95ef00c007ca852285efe02fb28a87a286130604043e899862a106a10793558700a38cb7fe93550701238db7fe93558701a38db7fe93550702238eb7fe93558702238ce7fea38eb7fe935507036193238fb7fea38fe7fee390c6fc7074ca852685ef00a00e4a8593050004efe02fab0145e6604664a66406692561828071c693f7f50f2300f5003307c500a30ff7fe894663fcc60aa300f5002301f500230ff7fea30ef7fe994663f1c60aa301f500230ef7fea14663fac60893f5f50f9b9785003307a0400d8bad9f198e9b950701ad9f2a97719a1cc3b305c70023aef5fe63f5c6065cc31cc723aaf5fe23acf5fee14663fcc604137847005cc71ccb5ccb1ccf6108939807029396070293d8080223a2f5fe23a4f5fe23a6f5fe23a8f5fe33060641fd474297c69663f0c7020116937706fe93870702ba9714e314e714eb14ef13070702e31af7fe8280397122fc26f84af44ef052ec56e85ae45ee093f735006387074069c2aa8719a06303062a83c60500850513f735002380d7007d1685076df793f637003e87cdea3d48637dc804930806ff6378180133e8b700137878006304083093d84800138f1800120f2e9f2e87be86832e0700032e4700032387000328c70023a0d60123a2c60123a4660023a606014107c106e31eeffc85089208c695c6973d8a137886001377460093762600058a630c080083a8050003a84500a107a10523ac17ff23ae07ff11c798419107910523aee7fe6391061e09c603c705002380e7006274c27422798279626ac26a226b826b216182807d476379c70a094883c805009841638806290d486386061d9306c6fe03c3150003c8250093f306ff13843700938435009382330123801701a38067002381070113d94600ae92a687a28803a8170083a5570083a697001b53870103a7d7009b1f88001b9f85009b9e86001b5888019bd585019bd686011b1e87003363f3013368e801b3e5d501b3e6c60123a0680023a2080123a4b80023a6d800c107c108e39657fa9307190092073516b385f40033067640a29793780601137886009376460013772600058a6384080883cb050003cb150083ca250003ca350083c9450003c9550083c4650003c4750083c3850083c2950083cfa50003cfb50083cec50003ced50003c3e50083c8f50023807701a380670123815701a381470123823701a382270123839700a383870023847700a38457002385f701a385e7012386d701a386c70123876700a3871701c105c1076304080483c2050083cf150003cf250083ce350003ce450003c3550083c8650003c8750023805700a380f7012381e701a381d7012382c701a382670023831701a3830701a105a1079dc203c3050083c8150003c8250083c6350023806700a380170123810701a381d70091059107e30307e283c6050003c715008907238fd7fea38fe7fe890539b513f73700e31d07ec39b59306c6fe93f306ff1384170093841500938213012380170113d94600ae92a687a28803a8370083a5770083a6b7001b53870003a7f7009b1f88011b9f85019b9e86011b5888009bd585009bd686001b1e87013363f3013368e801b3e5d501b3e6c60123a0680023a2080123a4b80023a6d800c107c108e39657fa9307190092073d16b385f40033067640a297a1b593d84800938e18002e88033e88000333080085062334c7012330670041084107e3e5d6ff85089208c695c6973d8a01bb9306c6fe03c8150093f306ff13842700938425009382230123801701a380070113d94600ae92a687a28803a8270083a5670083a6a7001b53070103a7e7009b1f08011b9f05019b9e06011b5808019bd505019bd606011b1e07013363f3013368e801b3e5d501b3e6c60123a0680023a2080123a4b80023a6d800c107c108e39657fa9307190092073916b385f40033067640a29749b3aa8709b919ca0347050083c705007d166317f700050585057df6014582800345050083c705001d9d8280aa862e87b287630db50cb388c5403308c040b388a84006082e832a8e6372181b3346b5001d8a637fb50a63010612cdcb1386f7ff9d4563f8c51813061700b305c54093b5750093c5150093f5f50f638a0516b365e5009d896395051693f587ffba95033603002103210e233ccefee39a65fe13f687ff13f57700aa87b385c600329739cd0345070005462380a5006389c704034517000946a380a5006382c704034527000d462381a500638bc702034537001146a381a5006384c7020345470015462382a500638dc700034557001946a382a5006386c700834767002383f5003685828029ea3306f5001d8a65ca1386f7fffdd7b307c5007d5821a07d16e30106ffb305c70003c5050093f57700fd17a380a700e5f59d4763fac70ab2871d48e117b305f7008861b385f60088e1e369f8fe93777600cdd7fd173306f700834506003386f6002300b600f5b71376750041ca9385f7ffc9d72a867d5821a0fd15e38005f903450700050693777600a30fa6fe0507edf79d4763fcb704938885ff93f888ffa10833051601ba8703b807002106a107233c06ffe31aa6fe469793f77500130617008ddfba9711a005060347f6ff0505a30fe5fee31af6fe36858280cdba3685d5b713061700f9bfb287a5b73285ae8713061700e1f919b73e8625bf2a86be8549bf000000000000cdccccccccccccccd182e6ad7f520e5108c9bcf367e6096a1f6c3e2b8c68059b3ba7ca8485ae67bb6bbd41fbabd9831f2bf894fe72f36e3c79217e1319cde05bf1361d5f3af54fa54b598638d6c56d340101010101010101ff00ff00ff00ff00fffefefefefefefe80808080808080800a0a0a0a0a0a0a0aaf47e17a14ae4701555555555555555533333333333333330f0f0f0f0f0f0f0f01010101010101019a9999999999990100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000a0da0a000000000000100000000000000400000000000000a0ca020000000000001008000000000040000000000000000100000000000000300a010000000000000000000000000030b2020000000000011101250e1305030e10171b0eb44219110155170000023901030e0000032e001101120640186e0e030e3a0b3b053f198701190000042e00110112064018030e3a0b3b05360b3f198701190000052e006e0e030e3a0b3b05200b0000062e001101120640186e0e030e3a0b3b050000072e006e0e030e3a0b3b0b200b0000082e011101120640186e0e030e3a0b3b0b360b0000091d00311311011206580b590b570b00000a1d0031135517580b590b570b00000b1d00311311011206580b5905570b00000c1d0031135517580b5905570b00000d2e006e0e030e3a0b3b0b3f19200b00000e2e011101120640186e0e030e3a0b3b0b3f1900000f1d0131135517580b590b570b0000101d01311311011206580b590b570b0000111d01311311011206580b5905570b0000121d0131135517580b5905570b0000132e006e0e030e3a0b3b053f19200b0000142e011101120640186e0e030e3a0b3b05360b3f190000152e011101120640186e0e030e3a0b3b053f190000162e0111011206401831130000172e0011011206401831130000182e001101120640186e0e030e3a0b3b0b0000192e011101120640186e0e030e3a0b3b0b00001a2e011101120640186e0e030e3a0b3b0500001b2e011101120640186e0e030e3a0b3b05360b3f1987011900001c2e001101120640186e0e030e3a0b3b0b3f1987011900001d2e006e0e030e3a0b3b0b870119200b00001e2e001101120640186e0e030e3a0b3b0b360b3f19870119000000700000000400000000000801752b00001c0060460000000000002b13000000000000000000007011000002742f0000020000000003326e0100000000000e00000001527c4f000064380000010b020002742f000002953f000004406e0100000000000e0000000152190f0000028e010300000000242600000400000000000801752b00001c005a170000880000002b1300000000000000000000a0110000023b1a00000284050000052f0d00009017000002f90501062eb3010000000000020000000152dc350000dd0c000002eb0102ab3f0000029733000005e6380000182500000593030105e6380000182500000593030105e6380000182500000593030105e6380000182500000593030105e63800001825000005930301059a2a00006c2300000593030105eb2c0000d14900000593030105ba3b00006f3a00000593030105770c0000f90300000536050105e638000018250000059303010000025f0d0000029733000005ae420000182500000701040105ae420000182500000701040105ae420000182500000701040105ae420000182500000701040105ae420000182500000701040105b03300008d1800000701040105ff0b0000d537000007010401000005a6000000794a00000273040105fd13000057440000027304010524490000900500000249050105b8080000cc00000002490501050b2a0000f903000002610601000293330000025b130000029034000007fd4b00005429000003d00100027b4100000736140000c8490000038e01078f3e000093330000038901078f3e000093330000038901000002544c0000024f3100000830b3010000000000420100000152fc1600007638000004d3030965000000a0b30100000000000200000004f1360ac61b00000000000004f1150972000000b2b30100000000000200000004f2360ad31b00004000000004f215097f000000fab30100000000000200000004fd360ae01b00007000000004fd1509f300000008b40100000000000200000004fd470b0001000022b4010000000000020000000403011e0b8c00000034b401000000000002000000040701360ced1b0000a0000000040701150b0d01000042b401000000000002000000040701470b1a01000050b401000000000006000000040f0133000002550c000007472d0000c03e000004430107441b0000f204000004430107c1160000b410000004430107aa3000004e2b000004430100022a2b00000d01150000581d000004870100028b4700000dc54a00001d3c0000042a010002761500000efebb010000000000700000000152ef30000093330000049a0fd902000020090000049b11103c1d000004bc01000000000008000000044e1d11a71c000004bc0100000000000800000019f80209094101000004bc010000000000080000001bef5000000a0f0300005009000004511c09ec21000016bc01000000000004000000045116092103000024bc010000000000080000000451280fd824000080090000046514120b1e0000b0090000225901090af81d0000e0090000171209000000000002c60700000d73350000581d000004870100020f0f00000ed6c2010000000000720000000152f528000093330000049a0fe5020000100e0000049b1110901d0000dcc201000000000008000000044e1d11a71c0000dcc20100000000000800000019f802090941010000dcc2010000000000080000001bef5000000afa030000400e000004511c09f9210000f2c20100000000000400000004511609b11b0000fec201000000000008000000044f190fe5240000700e000004651412171e0000a00e0000225901090af81d0000d00e00001712090000000000024b4800000e48c3010000000000720000000152af48000093330000049a0ff1020000000f0000049b11109d1d00004ec301000000000008000000044e1d11a71c00004ec30100000000000800000019f8020909410100004ec3010000000000080000001bef5000000a0f030000300f000004511c090622000064c30100000000000400000004511609b11b000070c301000000000008000000044f190ff2240000600f000004651412231e0000900f0000225901090af81d0000c00f0000171209000000000002210800000e72c40100000000007000000001521f03000093330000049a0ffd02000080100000049b1110aa1d000078c401000000000008000000044e1d11a71c000078c40100000000000800000019f80209094101000078c4010000000000080000001bef5000000afa030000b010000004511c09132200008ac401000000000004000000045116092103000098c4010000000000080000000451280fff240000e0100000046514122f1e000010110000225901090af81d00004011000017120900000000000002d74d000013e90a00001e0b000008bd0601137f0300005331000008f6060113c94c00004344000008100701056b0d000088050000086e05011472b4010000000000e4010000015289020000cc34000008de04030b6206000090b40100000000000c00000008e504130b6f060000acb40100000000000400000008ea04190b7c060000e8b401000000000002000000080a051a1289060000d00000000817052411df1f0000d0b5010000000000040000000880051211cc1f0000d0b5010000000000040000000ec702090b32220000d0b5010000000000020000000e6d020c000000121b13000010010000081a051112ec1f0000400100000894041212cc1f0000700100000ec702090c32220000a00100000e6d020c00000012c8210000d0010000080b05200b5001000062b501000000000006000000139403160b6a01000076b501000000000004000000139503090012d521000000020000080c05210b5d01000068b501000000000004000000139403160b770100007ab5010000000000040000001395030900118906000094b50100000000001a000000080e052411df1f00009ab5010000000000040000000880051211cc1f00009ab5010000000000040000000ec702090b322200009ab5010000000000040000000e6d020c0000001184200000beb40100000000001c00000008eb0416101f200000beb40100000000001c0000001231091013200000beb40100000000001c00000011200910771f0000beb40100000000001c00000011874c10ea1e0000beb40100000000001c000000105331111d1f0000beb40100000000001c0000000a940d09104d1f0000beb40100000000001c0000000c321110dd1e0000beb40100000000001c0000000f7c09120a1c0000300200000ab0091d104c1c0000cab401000000000002000000092b350927010000cab4010000000000020000000953520000125f1f0000800200000ab10915108d1f0000ccb4010000000000080000000f541c1030200000ccb40100000000000800000010501609db200000ccb40100000000000800000011871f0000092e1f0000d6b4010000000000020000000f54150000000000000000000015acb6010000000000780300000152784b0000e5300000083c0512a6220000b0020000083e05170c99220000e00200001483020f001136210000dab601000000000004000000084705251129210000dab6010000000000040000001641033311ba1c0000dab6010000000000040000001608032711581c0000dab60100000000000400000019e502090999000000dab6010000000000040000001b62500000000011041f0000deb6010000000000da0000000847052311f71e0000deb60100000000006e0000000a8b010912a2200000100300000a5801100f9020000040030000128c190fe720000070030000122c12090a1c000002b7010000000000040000000b260e09ff2000001ab7010000000000040000000b3212090b21000026b70100000000000a0000000b391309172100003cb70100000000000a0000000b412509f320000016b7010000000000040000000b2e1000000011f91f0000feb6010000000000040000000a57011211cc1f0000feb6010000000000040000000ec702090b32220000feb6010000000000020000000e6d020c00000011a22000006ab70100000000004e0000000a8c010910902000006ab70100000000004a000000128c1910e72000006ab70100000000004a000000122c12090a1c00006ab7010000000000040000000b260e0917210000a2b70100000000000c0000000b4125090b21000096b7010000000000040000000b391309ff20000092b7010000000000040000000b321200000000124f210000a0030000084c05131274210000d003000016b901091143210000b8b7010000000000120000001814010c10c71c0000beb70100000000000400000016dc1f0bc21d0000beb701000000000004000000195a010f000000000cb322000000040000084c051c1184200000ecb70100000000007201000008590523101f200000ecb7010000000000720100001231091013200000f2b70100000000001e00000011200910771f0000f2b70100000000001e00000011874c10ea1e0000f2b70100000000001e000000105331111d1f0000f2b70100000000001e0000000a940d09104d1f0000f2b70100000000001e0000000c321110dd1e0000f2b70100000000001e0000000f7c09120a1c0000300400000ab0091d104c1c0000feb701000000000002000000092b350927010000feb7010000000000020000000953520000125f1f0000800400000ab10915108d1f000000b8010000000000080000000f541c103020000000b80100000000000800000010501609db20000000b80100000000000800000011871f0000092e1f00000ab8010000000000020000000f541500000000000000103d20000010b80100000000004e01000011220910d41c000010b801000000000014000000113a270b8401000010b80100000000000600000019d60d1f11ee1c000016b80100000000000800000019da0d200be11c000016b80100000000000800000019460617000bfb1c00001eb80100000000000600000019db0d2400101320000024b80100000000001a00000011471510771f000024b80100000000001a00000011874c10ea1e000024b80100000000001a000000105331111d1f000024b80100000000001a0000000a940d09104d1f000024b80100000000001a0000000c321110dd1e000024b80100000000001a0000000f7c09120a1c0000b00400000ab0091d104c1c00002eb801000000000002000000092b3509270100002eb8010000000000020000000953520000125f1f0000000500000ab10915108d1f000030b8010000000000080000000f541c103020000030b80100000000000800000010501609db20000030b80100000000000800000011871f0000092e1f00003ab8010000000000020000000f541500000000000000101320000040b80100000000001c00000011473510771f000040b80100000000001c00000011874c10ea1e000040b80100000000001c000000105331111d1f000040b80100000000001c0000000a940d09104d1f000040b80100000000001c0000000c321110dd1e000040b80100000000001c0000000f7c09120a1c0000300500000ab0091d104c1c00004cb801000000000002000000092b3509270100004cb8010000000000020000000953520000125f1f0000800500000ab10915108d1f00004eb8010000000000080000000f541c10302000004eb80100000000000800000010501609db2000004eb80100000000000800000011871f0000092e1f000058b8010000000000020000000f541500000000000000104920000092b801000000000012000000115a12091f2300009eb801000000000004000000117f0e0010951c0000c0b80100000000000600000011501910151d0000c0b8010000000000060000001b1a0e11641c0000c0b80100000000000600000019e5020909a6000000c0b8010000000000060000001b62500000000a161c0000b00500001150190a55200000f005000011541b0f221c00006006000011631a10701c000032b901000000000002000000092b35093401000032b9010000000000020000000953520000096120000034b90100000000000c00000011641b106d2000004ab901000000000012000000116616092c23000056b901000000000004000000117f0e0009081d0000bcb801000000000004000000114f2c10821c0000a8b801000000000010000000114a121181220000b4b8010000000000040000001bcb051b1173220000b4b8010000000000040000000d7e04080b61220000b4b8010000000000040000000d2e03090000000000001289060000b00600000863052811df1f0000bab9010000000000040000000880051211cc1f0000bab9010000000000040000000ec702090b32220000bab9010000000000020000000e6d020c000000111b130000e6b9010000000000260000000865051512ec1f0000f00600000894041212cc1f0000200700000ec702090c32220000500700000e6d020c000000000d8b3b00000430000008f20113981800003d2d000008f4050113123400001d2b00000843070105c1280000ea1d0000089c04011630c20100000000009800000001520813000011ca1900003cc20100000000001800000008e6071b0b0b1200003cc20100000000000c0000001f17011200116718000062c20100000000005800000008e8070911ac2400006cc20100000000004a0000001f650127115b1700006ec20100000000004800000020270516116f17000082c2010000000000060000001f66013c0b6f06000082c2010000000000060000001f700109000b0b1200008ac2010000000000140000001f6701150b0b120000a0c2010000000000160000001f6901110000000013db070000fe24000008e507010002c51b00000559180000e7310000089304010002ed31000002cc3400000656b6010000000000560000000152874d00007f1b000008f304000005ac090000434d0000086404010517100000d1090000087904011532ba0100000000007e0100000152943c0000e73100000838040cff110000800700000839041912a71f0000b0070000084d041d0a2e1c0000e00700001d2f1100124f130000100800000856041a115c130000baba01000000000018000000086b04150bb3010000c0ba010000000000120000000881042c00115c130000e0ba01000000000018000000086c04190bb3010000e6ba010000000000120000000881042c0011221d000000bb010000000000040000000873041f11ce1d000000bb010000000000040000001996011a09b300000000bb0100000000000400000017ee1c00000bbf01000004bb010000000000080000000876040b0012b31f000040080000083f041d0a3a1c0000700800001d2f11000bcb01000052bb0100000000000a00000008460415122f1d0000a0080000085d042612da1d0000e0080000195a010f10e61d000080bb0100000000000400000017d93609c000000080bb0100000000000400000017ee1c0000000002f101000007244000000c3c00001f5501023b3b00000e6ebc010000000000bc01000001527e3800003d2d00001f1f0fc7200000100a00001f201212b4200000400a0000123f050911b3210000f4bc010000000000d40000001272020f11561d0000febc01000000000008000000249e01320b411e0000febc01000000000008000000195a010900118b1e000006bd010000000000ac00000024a2012209971e00000cbd0100000000001a000000252c1010a31e000026bd0100000000008c000000252f0510cd00000026bd0100000000000c0000002552160b8401000026bd0100000000000c000000054005160010bb1e00006cbd0100000000000a000000256a1609462300006cbd010000000000020000002514070010af1e000056bd0100000000000a000000256916093923000056bd010000000000020000002514070009da0000004abd0100000000000400000025651b09971e00009ebd0100000000001400000025771609971e00007ebd01000000000012000000255a1e000011631d0000bebd0100000000000200000024b701430b411e0000bebd01000000000002000000195a0109001152220000c0bd0100000000000400000024b8011c11781e0000c0bd010000000000040000000da9050d095a1e0000c0bd01000000000004000000231a0900000000000f5c210000700a00001f252712a0210000a00a0000165f040d128d210000d00a00002445022912491d0000000b000024de03091145220000d0bc0100000000000a00000019090913116c1e0000d0bc0100000000000a0000000da9050d095a1e0000d0bc0100000000000a000000231a09000000000000000002b140000002454800000592040000542900001f35010100023d1b000005a3240000542900001f650101000002432b000005474d0000664a00001f6f01011510c00100000000002001000001526f0a0000454800001f34011292240000b00b00001f350123114817000034c0010000000000de00000020270516126f170000e00b00001f3601100c6f060000100c00001f700109000b0b1200005cc0010000000000160000001f3801150c0b120000400c00001f4101110bbf24000092c0010000000000020000001f410111127a180000700c00001f3c01220f25120000b00c00001f1a091191180000b2c00100000000000a00000008a3041209c0220000b2c00100000000000a0000001f1a260000000b0b120000fec0010000000000120000001f3e011100000013641e00003d1b00001f63010100026d4b000007291e00000f3000001f15010002a3090000020f300000070b380000542900001f1a01000002321b00000514300000ec0400001f7b010105cf0e0000664a00001f9101010002114d000002ec0400000550300000542900001f7c0101000002dc3a00001530c10100000000000001000001524b050000ec0400001fd40112a4180000f00c00001fd50109129f240000200d00001f7c012311c91800006cc1010000000000c40000002027051612b1180000500d00001f7d01100c6f060000800d00001f920109000b0b12000080c1010000000000180000001f8801150b0b120000a6c1010000000000180000001f7f0115127a180000b00d00001f8301220f25120000e00d00001f1a091191180000d2c10100000000000a00000008a3041209c0220000d2c10100000000000a0000001f1a260000000b0b1200001ac2010000000000160000001f85011100000000000555340000932400001f1301010002d4320000162abe010000000000b400000001523c1a0000101626000038be0100000000009600000008a41a110426000038be010000000000960000002679022a0cf7250000300b000026b6060f00000017debe010000000000380000000152481a000007ae190000da32000008a3010714480000514f000008bf010002973300001816bf0100000000000a0000000152a74b00007745000008c61920bf010000000000b60000000152a2450000da32000008ca103c1a00002ebf010000000000a200000008cb09101626000030bf0100000000009600000008a41a110426000030bf010000000000960000002679022a0cf7250000700b000026b6060f0000000019d6bf0100000000003a0000000152e53a0000514f000008ce09481a0000f6bf0100000000001400000008cf090000022a0a000005da1000009333000008bb09010002d30c00001abac30100000000001600000001524b3300002511000008d0080b0e1b0000bac30100000000001600000008d0083e00000002db3c000002ce4d0000024d4c0000192ab3010000000000040000000152340a0000b54f000001fa10a10100002ab30100000000000400000001fa0509340000002ab30100000000000200000003d21e0000000002242f000002d0070000052a2f0000b01000002742020100000002df3c000005ab0a00008e110000065f0a0105ab0a00008e110000065f0a0105ab0a00008e110000065f0a0105ab0a00008e110000065f0a0100029d34000002a11e0000022025000007663600000e490000097c0107153e0000c1010000097c0107712c000076440000097c01076b4e00005a410000097c0107a01c000006400000097c010002383900000712000000a41b0000094b0107812f0000094d00001b5b0107e13400007c2300001b5b01078c2300004b370000094b010002614e000005ef390000764400001bc7050100029733000007740b0000ff3d00001b190100024d0c0000071a1d00002c4500001bd90100000297330000058a120000d11b000019e4020105501c0000fc2900001956010105404700009a4a000019cb0d01052c270000fb400000199806010518060000124100001942060105924400006209000019860d01053a2a0000862a00001916040105443b0000ee3d000019e4020105b41a0000d1120000198f010105e64400002f3200001956010105c6270000da09000019f70201055b0e00002b19000019040901054c0400000a1b000019560101054c0400000a1b00001956010102b607000003c8c20100000000000e0000000152fa450000c93c0000190b0d0005c6270000da09000019f7020105c6270000da09000019f7020105c6270000da09000019f702010002b4030000023b3b000007af050000d934000017d7010761370000f62a000017e30107f20d0000ff12000017d7010784410000fe33000017e3010002793a000005fa010000ee49000017ec01010002973300000740320000cd1800001711010740320000cd1800001711010740320000cd1800001711010740320000cd1800001711010002b140000005e9150000d9340000175f01010000029e0d000002114d00000780150000e73e0000235201000297330000075e1d0000a6400000231901075e1d0000a64000002319010000020830000007391900000830000025290107f53e00002d3f00002534010d2c4b0000db1d00002547010772100000f84100002513010772100000f8410000251301000002a11e0000027a2f000002b62b00000298460000055e1300002b2500000aaa090105b53f0000fc4200000a8f0d01057b390000f60000000a56010105ec080000b60f00000a8a0101000002a611000002ac1100000760290000ea3c00000c310102670d000007cf430000b61100000c35010000000002704a0000025d310000023b3b00000761310000a61e00000f78010002e84d000007ad460000c32000000f5401000002e14d0000023b3b0000072b0800009e130000104d01020c000000021749000007a5170000590000001050010000000002961c000002a30900000763060000822700001d2e01076c140000d32300001d2e0100000002df080000023b3b0000054b490000712200000e6c02010002844a00000582220000764400000ec602010582220000764400000ec602010582220000764400000ec602010000000208000000020c0000000d280b00008c1b000011860107230f0000a1460000111a01028c1b0000076520000054290000118701000d2b090000a51a0000112601071f41000023140000117a01072a2c0000d2010000117201072a2c0000d2010000117201071f41000023140000117a010002a11e0000029733000007584c00000c00000012300107f14d00001f0100001229010002114d000007da1b00001f010000128a010002bb3200000517280000620c0000126c020100025a45000005e82d0000c9320000123e0501000002680b000007ba400000f43f00000b180107bf2b0000c23900000b240107d80f0000fe2b00000b0b010717230000592300000b11010717230000592300000b11010717230000592300000b1101000297330000053d390000e33600001607030105b62900008d4a00001640030107a80d00000e2c000016d30105e93600002537000016b80101050a04000096400000165b040100027a2f000002a73300000524010000ab05000018130101000002174b0000022a2b000005e54e00001f4b000024dd03010002844a000005652800001f4b000024410201000297330000056a2e000026350000249b0101000000022049000005b63d0000b71b0000138f030105a3340000570f0000138f030102822d0000026a15000005bd470000bb4a000021e8010105bd470000bb4a000021e8010105bd470000bb4a000021e8010105bd470000bb4a000021e80101000000029e0d000002a20d000002ec00000005401a0000e03600000d53050100028a24000005233c0000342b00000da8050105233c0000342b00000da8050100000595470000f63100000d930401026b3a0000051a4d00001f2c00000d2a030100057e0900001f2c00000d7d04010002e508000002a033000005790f00009c050000145602010503470000df3d00001482020105ba0300008244000014bb030105f6060000a70e000014120601001be2bb0100000000000e00000001527b420000bb3c0000148b0703117f230000e4bb0100000000000c000000148c07050973230000e4bb0100000000000c0000001c860500000002544c0000028b47000005bc2f0000ae4a00001ae4040105bc2f0000ae4a00001ae40401051e4a0000444f00001acd0401051e4a0000444f00001acd0401000002ec2a00001c24ba0100000000000e00000001522d170000e93000001c6e1d60400000091300001c95011d411000004b3400001c85011ef0bb0100000000000e000000015210330000644500001c50030002051b000002bc27000015b0bb01000000000012000000015255480000933300001ebb021118120000b0bb010000000000120000001ebc021b11dd140000b0bb0100000000001200000008440709090b120000b0bb010000000000120000001f591200000000021c35000015c2bb010000000000120000000152c2020000933300001ed6021118120000c2bb010000000000120000001ed7021b11dd140000c2bb0100000000001200000008440709090b120000c2bb010000000000120000001f5912000000000002fa14000003d4bb0100000000000e0000000152180500001d13000020720602664b00000531350000e1190000202505010532070000823a00002025050105740700003a3f000020250501000206330000050b4200000d0a0000209b0701000002112800000221190000050a2400008f2d000022580101050a2400008f2d000022580101050a2400008f2d000022580101050a2400008f2d0000225801010002063300000ed0c3010000000000a200000001522d1100009333000022830f08130000f00f000022830a12ca1900002010000008e6071b0c0b120000501000001f1701120011671800000ec40100000000005800000008e8070911ac24000018c40100000000004a0000001f650127115b1700001ac40100000000004800000020270516116f1700002ec4010000000000060000001f66013c0b6f0600002ec4010000000000060000001f700109000b0b12000036c4010000000000140000001f6701150b0b1200004cc4010000000000160000001f6901110000000000000002f1060000020338000005e12e00006a190000269906010573190000142f000026b5060102973300000572160000084800002677020100000000003c0000000200000000000800ffffffff326e0100000000000e00000000000000406e0100000000000e0000000000000000000000000000000000000000000000ec0100000200740000000800ffffffff2ab301000000000004000000000000002eb3010000000000020000000000000030b3010000000000420100000000000072b4010000000000e40100000000000056b60100000000005600000000000000acb6010000000000780300000000000024ba0100000000000e0000000000000032ba0100000000007e01000000000000b0bb0100000000001200000000000000c2bb0100000000001200000000000000d4bb0100000000000e00000000000000e2bb0100000000000e00000000000000f0bb0100000000000e00000000000000febb01000000000070000000000000006ebc010000000000bc010000000000002abe010000000000b400000000000000debe010000000000380000000000000016bf0100000000000a0000000000000020bf010000000000b600000000000000d6bf0100000000003a0000000000000010c0010000000000200100000000000030c1010000000000000100000000000030c20100000000009800000000000000c8c20100000000000e00000000000000d6c2010000000000720000000000000048c30100000000007200000000000000bac30100000000001600000000000000d0c3010000000000a20000000000000072c4010000000000700000000000000000000000000000000000000000000000a2b3010000000000a6b3010000000000aab3010000000000b2b3010000000000beb3010000000000c2b301000000000000000000000000000000000000000000b4b3010000000000bcb3010000000000c2b3010000000000cab301000000000000000000000000000000000000000000fcb301000000000008b40100000000000ab401000000000014b40100000000000000000000000000000000000000000036b401000000000042b401000000000044b40100000000004cb401000000000000000000000000000000000000000000ecb4010000000000f2b4010000000000f6b4010000000000fcb4010000000000b0b5010000000000e0b50100000000000000000000000000000000000000000010b601000000000030b601000000000050b601000000000056b60100000000000000000000000000000000000000000018b601000000000020b601000000000050b601000000000056b60100000000000000000000000000000000000000000018b601000000000020b601000000000050b601000000000056b60100000000000000000000000000000000000000000018b601000000000020b601000000000050b601000000000056b60100000000000000000000000000000000000000000062b501000000000068b501000000000076b50100000000007ab50100000000000000000000000000000000000000000068b50100000000006cb50100000000007ab50100000000007eb501000000000000000000000000000000000000000000beb4010000000000c2b4010000000000cab4010000000000ccb4010000000000d4b4010000000000d6b4010000000000d8b4010000000000dab401000000000000000000000000000000000000000000ccb4010000000000d4b4010000000000d6b4010000000000d8b401000000000000000000000000000000000000000000aeb6010000000000c4b6010000000000c6b6010000000000ceb601000000000000000000000000000000000000000000aeb6010000000000c4b6010000000000c6b6010000000000ceb601000000000000000000000000000000000000000000f0b6010000000000fab601000000000002b70100000000004cb701000000000000000000000000000000000000000000f0b6010000000000f4b601000000000002b701000000000048b701000000000000000000000000000000000000000000f0b6010000000000f4b601000000000002b701000000000048b701000000000000000000000000000000000000000000b8b7010000000000ceb7010000000000d4b7010000000000d8b701000000000000000000000000000000000000000000b8b7010000000000ceb7010000000000d4b7010000000000d8b701000000000000000000000000000000000000000000d0b7010000000000d4b7010000000000dab7010000000000dcb701000000000000000000000000000000000000000000f2b7010000000000f6b7010000000000feb701000000000000b801000000000008b80100000000000ab80100000000000cb801000000000010b80100000000000000000000000000000000000000000000b801000000000008b80100000000000ab80100000000000cb80100000000000000000000000000000000000000000024b801000000000028b80100000000002eb801000000000030b801000000000038b80100000000003ab80100000000003cb80100000000003eb80100000000000000000000000000000000000000000030b801000000000038b80100000000003ab80100000000003cb80100000000000000000000000000000000000000000040b801000000000042b80100000000004cb80100000000004eb801000000000056b801000000000058b80100000000005ab80100000000005cb8010000000000000000000000000000000000000000004eb801000000000056b801000000000058b80100000000005ab801000000000000000000000000000000000000000000c6b8010000000000c8b80100000000000cb901000000000010b901000000000012b901000000000018b901000000000000000000000000000000000000000000d0b8010000000000d8b8010000000000dab8010000000000deb8010000000000e0b8010000000000e6b8010000000000e8b8010000000000f8b8010000000000fab8010000000000fcb801000000000000b90100000000000cb90100000000000000000000000000000000000000000018b901000000000030b901000000000032b901000000000034b901000000000040b901000000000042b901000000000044b901000000000048b90100000000000000000000000000000000000000000062b901000000000068b90100000000006cb901000000000072b901000000000098b9010000000000cab901000000000000000000000000000000000000000000eeb9010000000000f6b901000000000008ba0100000000000cba01000000000000000000000000000000000000000000eeb9010000000000f6b901000000000008ba0100000000000cba01000000000000000000000000000000000000000000eeb9010000000000f2b901000000000008ba0100000000000cba010000000000000000000000000000000000000000004aba01000000000052ba01000000000056ba0100000000005eba0100000000000000000000000000000000000000000064ba0100000000008eba0100000000000ebb0100000000001ebb0100000000000000000000000000000000000000000064ba0100000000008eba0100000000000ebb0100000000001ebb01000000000000000000000000000000000000000000a0ba010000000000aeba010000000000b2ba0100000000000cbb0100000000000000000000000000000000000000000022bb01000000000040bb0100000000005ebb01000000000068bb0100000000000000000000000000000000000000000022bb01000000000040bb0100000000005ebb01000000000068bb010000000000000000000000000000000000000000006cbb01000000000072bb01000000000078bb0100000000007cbb01000000000080bb01000000000084bb010000000000000000000000000000000000000000006cbb01000000000072bb01000000000078bb0100000000007cbb01000000000080bb01000000000084bb0100000000000000000000000000000000000000000004bc0100000000005abc01000000000060bc0100000000006ebc0100000000000000000000000000000000000000000014bc01000000000016bc0100000000002cbc01000000000030bc010000000000000000000000000000000000000000003abc01000000000044bc01000000000060bc0100000000006ebc010000000000000000000000000000000000000000003abc01000000000044bc01000000000060bc0100000000006ebc010000000000000000000000000000000000000000003abc01000000000044bc01000000000060bc0100000000006ebc01000000000000000000000000000000000000000000b4bc010000000000ccbc010000000000ecbc010000000000c8bd01000000000000000000000000000000000000000000b4bc010000000000ccbc010000000000ecbc010000000000c8bd01000000000000000000000000000000000000000000ccbc010000000000dabc010000000000f8bd010000000000fcbd01000000000000000000000000000000000000000000ccbc010000000000dabc010000000000f8bd010000000000fcbd01000000000000000000000000000000000000000000ccbc010000000000dabc010000000000f8bd010000000000fcbd01000000000000000000000000000000000000000000ccbc010000000000dabc010000000000f8bd010000000000fcbd0100000000000000000000000000000000000000000038be0100000000003cbe01000000000044be0100000000004abe01000000000066be0100000000006cbe0100000000000000000000000000000000000000000030bf01000000000034bf0100000000003cbf01000000000042bf0100000000005ebf01000000000064bf0100000000000000000000000000000000000000000026c001000000000028c001000000000034c001000000000012c10100000000000000000000000000000000000000000038c00100000000003cc001000000000040c001000000000044c00100000000000000000000000000000000000000000038c00100000000003cc001000000000040c001000000000044c00100000000000000000000000000000000000000000082c00100000000008cc00100000000008ec001000000000092c001000000000000000000000000000000000000000000a0c0010000000000a4c0010000000000aac0010000000000e8c0010000000000ecc0010000000000f6c001000000000000000000000000000000000000000000a0c0010000000000a4c0010000000000aac0010000000000e8c0010000000000ecc0010000000000f6c00100000000000000000000000000000000000000000042c101000000000054c10100000000006cc101000000000030c2010000000000000000000000000000000000000000004ac10100000000004cc10100000000006cc101000000000030c20100000000000000000000000000000000000000000070c101000000000074c101000000000078c10100000000007cc10100000000000000000000000000000000000000000070c101000000000074c101000000000078c10100000000007cc101000000000000000000000000000000000000000000c0c1010000000000c4c1010000000000cac101000000000012c201000000000000000000000000000000000000000000c0c1010000000000c4c1010000000000cac101000000000012c201000000000000000000000000000000000000000000dcc201000000000034c30100000000003ac301000000000048c301000000000000000000000000000000000000000000f0c2010000000000f2c201000000000006c30100000000000ac30100000000000000000000000000000000000000000014c30100000000001ec30100000000003ac301000000000048c30100000000000000000000000000000000000000000014c30100000000001ec30100000000003ac301000000000048c30100000000000000000000000000000000000000000014c30100000000001ec30100000000003ac301000000000048c3010000000000000000000000000000000000000000004ec3010000000000a6c3010000000000acc3010000000000bac30100000000000000000000000000000000000000000062c301000000000064c301000000000078c30100000000007cc30100000000000000000000000000000000000000000086c301000000000090c3010000000000acc3010000000000bac30100000000000000000000000000000000000000000086c301000000000090c3010000000000acc3010000000000bac30100000000000000000000000000000000000000000086c301000000000090c3010000000000acc3010000000000bac301000000000000000000000000000000000000000000dac3010000000000dcc3010000000000dec301000000000066c401000000000000000000000000000000000000000000dac3010000000000dcc3010000000000dec3010000000000fac301000000000000000000000000000000000000000000dac3010000000000dcc3010000000000dec3010000000000eec30100000000000000000000000000000000000000000078c4010000000000cec4010000000000d4c4010000000000e2c40100000000000000000000000000000000000000000088c40100000000008ac4010000000000a0c4010000000000a4c401000000000000000000000000000000000000000000aec4010000000000b8c4010000000000d4c4010000000000e2c401000000000000000000000000000000000000000000aec4010000000000b8c4010000000000d4c4010000000000e2c401000000000000000000000000000000000000000000aec4010000000000b8c4010000000000d4c4010000000000e2c401000000000000000000000000000000000000000000326e010000000000406e010000000000406e0100000000004e6e010000000000000000000000000000000000000000002ab30100000000002eb30100000000002eb301000000000030b301000000000030b301000000000072b401000000000072b401000000000056b601000000000056b6010000000000acb6010000000000acb601000000000024ba01000000000024ba01000000000032ba01000000000032ba010000000000b0bb010000000000b0bb010000000000c2bb010000000000c2bb010000000000d4bb010000000000d4bb010000000000e2bb010000000000e2bb010000000000f0bb010000000000f0bb010000000000febb010000000000febb0100000000006ebc0100000000006ebc0100000000002abe0100000000002abe010000000000debe010000000000debe01000000000016bf01000000000016bf01000000000020bf01000000000020bf010000000000d6bf010000000000d6bf01000000000010c001000000000010c001000000000030c101000000000030c101000000000030c201000000000030c2010000000000c8c2010000000000c8c2010000000000d6c2010000000000d6c201000000000048c301000000000048c3010000000000bac3010000000000bac3010000000000d0c3010000000000d0c301000000000072c401000000000072c4010000000000e2c4010000000000000000000000000000000000000000007261775f7665630073747200636f756e74005f5a4e34636f726535736c6963653469746572313349746572244c542454244754243134706f73745f696e635f73746172743137683231633736663939343638653065646545007b636c6f7375726523307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e005f5a4e34636f726533707472347265616431376831626239643039646638396234373532450077726974653c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e007b696d706c2335347d00616476616e63655f62793c636f72653a3a7374723a3a697465723a3a43686172496e64696365733e006e657874005f5a4e34636f726533737472367472616974733131305f244c5424696d706c2475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c5424737472244754242475323024666f722475323024636f72652e2e6f70732e2e72616e67652e2e52616e6765546f244c54247573697a652447542424475424336765743137683633326532303137643665353735396645006e6578743c5b7573697a653b20345d3e00636f6e7461696e735f6e6f6e5f636f6e74696e756174696f6e5f62797465006275696c64657273005f5a4e3131305f244c5424636f72652e2e6f70732e2e72616e67652e2e52616e676546726f6d244c54247573697a6524475424247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c54242475356224542475356424244754242447542435696e6465783137686163396536316662616530626263376145005f5a4e34636f726533666d7439466f726d617474657231327061645f696e74656772616c3137686238656639343965396131613633346545005f5a4e36335f244c5424636f72652e2e63656c6c2e2e426f72726f774d75744572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683636336332373865383138373636393045005f5a4e34636f726533666d74336e756d35335f244c5424696d706c2475323024636f72652e2e666d742e2e55707065724865782475323024666f7224753230246936342447542433666d743137683464336136353331313038303933376445005f5a4e34636f726533666d7439466f726d617474657239616c7465726e617465313768333537326537646636323036356664374500696e646578005f5a4e34636f7265366f7074696f6e31354f7074696f6e244c5424542447542439756e777261705f6f72313768343165333439646137383638346138334500616c69676e5f6f66667365743c75383e005f5a4e34636f72653373747232315f244c5424696d706c24753230247374722447542439656e64735f776974683137683139626662313333653233336465306145005f5a4e34636f726535736c69636532395f244c5424696d706c2475323024247535622454247535642424475424336765743137683233646638653962656438656665346645005f5a4e34636f726533666d74386275696c64657273313044656275675475706c65356669656c6432385f24753762242475376224636c6f7375726524753764242475376424313768636364396362623165623562613563364500656e74727900666d745f696e743c636f72653a3a666d743a3a6e756d3a3a55707065724865782c2075383e005f5a4e34636f726536726573756c743133756e777261705f6661696c65643137683030653934303161326339653536633045005f5a4e34636f726533666d74386275696c6465727338446562756753657435656e7472793137686531623638303262326163636539656445007074720070616464696e670077726974653c636861723e0069735f736f6d653c7573697a653e00676574005f5a4e37355f244c54247573697a65247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c542424753562245424753564242447542424475424336765743137683362336666656535366439303731313345005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243873706c69745f61743137683461343239666364306233623563343945005f5a4e3131305f244c5424636f72652e2e697465722e2e61646170746572732e2e656e756d65726174652e2e456e756d6572617465244c54244924475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e65787431376831623734616564656639323065303665450063686172005f5a4e34636f7265366f7074696f6e31354f7074696f6e244c5424542447542436696e736572743137686265366237313331636461646331646245005f5a4e34636f726536726573756c743139526573756c74244c542454244324452447542438616e645f7468656e3137683138643933303364393238646565393245005f5a4e34636f726536726573756c743139526573756c74244c542454244324452447542438616e645f7468656e313768316532623263316238653933626561654500636f70795f66726f6d5f736c696365007b696d706c2332397d007b696d706c233232357d005f5a4e34636f726533666d7439466f726d6174746572323564656275675f7475706c655f6669656c64315f66696e6973683137683963326264643732306464613133376545007b696d706c2336357d005f5a4e3130385f244c5424636f72652e2e697465722e2e61646170746572732e2e66696c7465722e2e46696c746572244c5424492443245024475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722447542435636f756e743137683631323362313132363938303130326445005f5a4e34636f72653370747235777269746531376830336462313664353065636536366165450072616e6765006f7074696f6e005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f72336e74683137683635613666633036633265613031396645005f5a4e34636f72653373747235636f756e743134646f5f636f756e745f6368617273313768653066306166323562653730356463664500616c69676e5f746f5f6f6666736574733c75382c207573697a653e005f5a4e34636f726533636d70336d696e3137683961303232643031326665326338333745007b696d706c23317d005f5a4e34636f726533666d743372756e313768666639613633333362396633663061614500676574636f756e7400697465725f6d75743c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e006272616e63683c28292c20636f72653a3a666d743a3a4572726f723e007b696d706c2332357d005f5a4e34636f7265336f70733866756e6374696f6e36466e4f6e63653963616c6c5f6f6e63653137683331326365396462383432326365623645005f5a4e34636f726533666d74386275696c64657273313044656275675475706c65356669656c643137686134393061356537663734366534656245005f5a4e34636f72653130696e7472696e736963733139636f70795f6e6f6e6f7665726c617070696e673137683165326664363834393232323263326345005f5a4e34636f726533666d7439466f726d6174746572397369676e5f706c75733137683765363563323535316433616561343445007369676e5f706c7573005f5a4e34636f72653373747235636f756e743233636861725f636f756e745f67656e6572616c5f6361736531376864313333363866323830386530613030450076616c69646174696f6e73005f5a4e34636f726535736c696365346974657238375f244c5424696d706c2475323024636f72652e2e697465722e2e7472616974732e2e636f6c6c6563742e2e496e746f4974657261746f722475323024666f7224753230242452462424753562245424753564242447542439696e746f5f697465723137683765326332623733366531386264656545005f5a4e34636f726533707472376d75745f70747233315f244c5424696d706c2475323024244250246d75742475323024542447542433616464313768333939313037663564323335643062374500497465724d75740047656e657269635261646978006e6578745f696e636c75736976653c636861723e005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243132616c69676e5f6f66667365743137686265366661383332613635626436303545007b696d706c2335337d0064726f705f696e5f706c6163653c26636f72653a3a697465723a3a61646170746572733a3a636f706965643a3a436f706965643c636f72653a3a736c6963653a3a697465723a3a497465723c75383e3e3e005f5a4e34636f7265337074723133726561645f766f6c6174696c653137683034656338646164326362346562306245006d75745f7074720073756d005f5a4e34636f726533666d7439466f726d61747465723770616464696e67313768386664646163386139653836623737364500636d7000696d706c73005f5a4e34636f72653373747232315f244c5424696d706c247532302473747224475424313669735f636861725f626f756e646172793137683034353265303532643135616334353245005f5a4e37355f244c54247573697a65247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c542424753562245424753564242447542424475424336765743137686337356165633633323166633531643545005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542439656e64735f77697468313768383363653331633938643238356662364500696e736572743c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e005f5a4e34636f726533666d74386275696c6465727331304465627567496e6e65723969735f7072657474793137683430666266303734623763353466303545007b696d706c2334317d005f5f72646c5f6f6f6d005f5a4e34636f72653373747235636f756e743131636f756e745f63686172733137683362393037393633646461313835376345007265706c6163653c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e005f5a4e34636f7265366f7074696f6e31354f7074696f6e244c542454244754243769735f736f6d653137686166353061376333383437653666373645006e74683c636f72653a3a7374723a3a697465723a3a43686172496e64696365733e005f5a4e34636f726533737472313176616c69646174696f6e733135757466385f66697273745f627974653137683962396637633933306431356335663945005f5a4e34636f726533666d7438676574636f756e743137683639663830313763343363306364653245005f5a4e34636f72653970616e69636b696e673970616e69635f7374723137683666303932373830653338346562353045005f5a4e34636f726535736c696365366d656d6368723138636f6e7461696e735f7a65726f5f6279746531376861303536386565313833303061353732450072656d00666d745f696e743c636f72653a3a666d743a3a6e756d3a3a4c6f7765724865782c2075383e005f5a4e34355f244c5424244c502424525024247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d74313768613430323766643039663261636331324500666d743c28293e005f5a4e36375f244c5424636f72652e2e61727261792e2e54727946726f6d536c6963654572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d74313768353264643636336235383463633535664500636f70795f6e6f6e6f7665726c617070696e673c75383e00616363756d007b696d706c2334387d007b636c6f7375726523307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542434697465723137686266616536663139613561623764656445006765745f756e636865636b65643c636f72653a3a666d743a3a72743a3a417267756d656e742c207573697a653e006765743c267374723e0070616e69635f646973706c61793c267374723e00756e777261705f6661696c6564002f72757374632f32663662633564323539653761623235646466646433336465353362383932373730323138393138007274005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f7234666f6c64313768623061333862663336373733633236364500636f756e743c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e005f5a4e34636f726533707472347265616431376831653634383335653639376533366630450073756d5f62797465735f696e5f7573697a65005f5a4e34636f726533666d7432727438417267756d656e743861735f7573697a653137686437613231613332353662616362386245005f5a4e3131305f244c5424636f72652e2e697465722e2e61646170746572732e2e656e756d65726174652e2e456e756d6572617465244c54244924475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e657874313768633030313137313163643937383139624500726573756c74005f5a4e37335f244c5424636f72652e2e666d742e2e6e756d2e2e4c6f776572486578247532302461732475323024636f72652e2e666d742e2e6e756d2e2e47656e657269635261646978244754243564696769743137686634306237613733623764393162653445004d61796265556e696e6974007b696d706c2336347d005f5a4e37335f244c54242475356224412475356424247532302461732475323024636f72652e2e736c6963652e2e636d702e2e536c6963655061727469616c4571244c542442244754242447542435657175616c3137686637383434376536346661643333376145005f5a4e3130365f244c5424636f72652e2e6f70732e2e72616e67652e2e52616e6765244c54247573697a6524475424247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c542424753562245424753564242447542424475424336765743137683761383664333261616263343034303345005f5a4e34636f72653463686172376d6574686f647332325f244c5424696d706c247532302463686172244754243131656e636f64655f757466383137683661333732316366346263313738623645005f5a4e34636f726533666d74336e756d313247656e65726963526164697837666d745f696e743137686363663535643038613665313532386645005f5a4e34636f726533666d74336e756d33696d7037666d745f7536343137683238366534643532373433386334363745005f5a4e34636f72653970616e69636b696e673570616e69633137686437373538656430613265383739363145006c6962726172792f636f72652f7372632f6c69622e72732f402f636f72652e353431663036343835316338633866372d6367752e3000726561645f766f6c6174696c653c7573697a653e005f5a4e3130385f244c5424636f72652e2e697465722e2e61646170746572732e2e66696c7465722e2e46696c746572244c5424492443245024475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722447542435636f756e7438746f5f7573697a6532385f24753762242475376224636c6f73757265247537642424753764243137686532646263323632336436376436643345005f5a4e34636f726533666d743131506f737450616464696e673577726974653137683130373832303864313037663934393045006164643c7573697a653e005f5a4e34636f726533666d7439466f726d61747465723977726974655f737472313768353330393765363135313339346565644500696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e2c20636f72653a3a6f70733a3a72616e67653a3a52616e676546726f6d3c7573697a653e3e007b696d706c2331357d00656e64735f776974683c75383e005f5a4e34636f726535736c696365366d656d636872366d656d6368723137683838333063653264646237323666636245006c656e5f75746638005f5a4e34636f72653463686172376d6574686f64733135656e636f64655f757466385f7261773137686230336466376165346464366562316445005f5a4e34636f726533666d74355772697465313077726974655f63686172313768666466623438666364333637346132384500616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23347d3a3a6669656c643a3a7b636c6f737572655f656e7623307d3e00636f7265005f5a4e34636f726533636d7035696d706c7335375f244c5424696d706c2475323024636f72652e2e636d702e2e5061727469616c4f72642475323024666f7224753230247573697a6524475424326c74313768383563303932356636663163316566654500646f5f636f756e745f6368617273005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542431336765745f756e636865636b656431376838333832313033623533356331333034450063656c6c006765743c75382c20636f72653a3a6f70733a3a72616e67653a3a52616e67653c7573697a653e3e004465627567496e6e65720066696e697368005f5a4e34636f726533666d74336e756d313247656e65726963526164697837666d745f696e7431376835383366363662653034373931303631450077726974655f70726566697800636861725f636f756e745f67656e6572616c5f6361736500706f73745f696e635f73746172743c75383e007265706c6163653c636861723e00506f737450616464696e6700697465723c75383e005f5a4e38375f244c5424636f72652e2e7374722e2e697465722e2e43686172496e6469636573247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683862646365633661316137393933386345005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542433676574313768396431656137353833353464396166364500656e756d6572617465005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683563636236663439653430616432356245005f5a4e34636f726535736c69636534697465723136497465724d7574244c54245424475424336e65773137683131393134666634646337396132326545006469676974005f5a4e34636f726535736c69636533636d7038315f244c5424696d706c2475323024636f72652e2e636d702e2e5061727469616c4571244c54242475356224422475356424244754242475323024666f7224753230242475356224412475356424244754243265713137683331383339323064643563373930336445006d656d6368725f616c69676e656400777261705f6275663c636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23317d3a3a777261703a3a7b636c6f737572655f656e7623307d3e005f5a4e34636f726533666d74386275696c6465727331305061644164617074657234777261703137686630613261643433323636313138356545005f5a4e34636f726533666d74386275696c64657273313044656275675475706c653666696e6973683137683262326465366164386361323965353845006974657200666f6c643c7573697a652c20636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c207573697a652c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e005f5a4e34636f72653373747235636f756e743233636861725f636f756e745f67656e6572616c5f6361736532385f24753762242475376224636c6f73757265247537642424753764243137686238333838383631636166343538396545007b636c6f7375726523307d3c2675382c207573697a652c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e00737065635f6e6578743c7573697a653e005f5a4e34636f726534697465723572616e67653130315f244c5424696d706c2475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722475323024666f722475323024636f72652e2e6f70732e2e72616e67652e2e52616e6765244c5424412447542424475424346e6578743137683166316635393732633862353338396245005f5a4e34636f726533737472313176616c69646174696f6e733138757466385f6163635f636f6e745f62797465313768386431353839303565613233346333334500757466385f6163635f636f6e745f62797465006164643c5b7573697a653b20345d3e006e65773c5b7573697a653b20345d3e005f5a4e34636f726535736c6963653469746572313349746572244c542454244754243134706f73745f696e635f73746172743137686632323465323937613136633263656145006e6578743c636f72653a3a736c6963653a3a697465723a3a497465723c636f72653a3a666d743a3a72743a3a417267756d656e743e3e005f5a4e34636f726535617272617938355f244c5424696d706c2475323024636f72652e2e6f70732e2e696e6465782e2e496e646578244c542449244754242475323024666f722475323024247535622454247533622424753230244e24753564242447542435696e6465783137683663646534633833393961376530333445007b696d706c23397d0064656275675f7475706c655f6e6577005f5a4e34636f726533666d74386275696c64657273313044656275675475706c653666696e69736832385f24753762242475376224636c6f737572652475376424247537642431376861393666623161373161643166373535450064656275675f7475706c655f6669656c64315f66696e697368006164643c75383e007b696d706c233138317d00666f6c643c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a6d61703a3a6d61705f666f6c643a3a7b636c6f737572655f656e7623307d3c2675382c207573697a652c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e3e005f5a4e34636f726535736c69636532395f244c5424696d706c2475323024247535622454247535642424475424313873706c69745f61745f756e636865636b65643137683765396534313435376636393734393145006e6578743c636f72653a3a736c6963653a3a697465723a3a497465723c636f72653a3a666d743a3a72743a3a506c616365686f6c6465723e3e007b696d706c2331377d005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542438697465725f6d75743137683030376635633136366631613761373245006172726179005f5a4e34636f7265337374723469746572323253706c6974496e7465726e616c244c5424502447542431346e6578745f696e636c75736976653137683938613230353930343932666138366445005f5a4e35325f244c542463686172247532302461732475323024636f72652e2e7374722e2e7061747465726e2e2e5061747465726e24475424313269735f7375666669785f6f663137683866653837336364343736333664316445005f5a4e34636f726533666d7439466f726d617474657238777261705f6275663137686636336162363038633262616362303045005f5a4e34636f726533666d74336e756d35325f244c5424696d706c2475323024636f72652e2e666d742e2e55707065724865782475323024666f72247532302469382447542433666d743137683438643832613435336137306166353745007b636c6f7375726523307d005f5a4e35365f244c54247573697a65247532302461732475323024636f72652e2e697465722e2e7472616974732e2e616363756d2e2e53756d244754243373756d3137683739356164323965353439386433333445005f5a4e34636f72653373747232315f244c5424696d706c2475323024737472244754243132636861725f696e64696365733137686466343535663065643137623532303045006765743c75382c207573697a653e005f5a4e34636f7265337074723132616c69676e5f6f66667365743137683534623332333739346162326331313545005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243961735f6368756e6b7331376831643562356538303063366463326238450061735f6368756e6b733c7573697a652c20343e005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243361646431376835666664656536393830656665666331450070616e69636b696e67006765745f756e636865636b65643c636f72653a3a666d743a3a72743a3a417267756d656e743e0064656275675f737472756374007b696d706c2332387d0065713c5b75385d2c205b75385d3e0044656275675475706c6500666d745f696e743c636f72653a3a666d743a3a6e756d3a3a55707065724865782c207536343e00636c616e67204c4c564d202872757374632076657273696f6e20312e37312e302d6e696768746c79202832663662633564323520323032332d30352d30392929006974657261746f72005f5a4e34636f726533737472313176616c69646174696f6e7331356e6578745f636f64655f706f696e74313768656364656330303032323838613566354500757466385f66697273745f627974650069735f636861725f626f756e64617279006d696e3c7573697a653e005f5a4e34636f72653373747235636f756e743330636f6e7461696e735f6e6f6e5f636f6e74696e756174696f6e5f627974653137686530636638653465356130663030393045005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137686134633765313364663063343439373145005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243361646431376833356564316564666234363437623138450077726974655f737472005f5a4e34636f726533666d74336e756d313247656e65726963526164697837666d745f696e743137686162643431393537653230363731373445006d617962655f756e696e697400696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e2c20636f72653a3a6f70733a3a72616e67653a3a52616e676546726f6d3c7573697a653e2c203132383e005f5a4e39395f244c5424636f72652e2e7374722e2e697465722e2e53706c6974496e636c7573697665244c54245024475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683536356238663563313134366339666645005f5a4e38315f244c5424636f72652e2e7374722e2e7061747465726e2e2e436861725365617263686572247532302461732475323024636f72652e2e7374722e2e7061747465726e2e2e53656172636865722447542431306e6578745f6d617463683137686231353436643361613035653433333145005f5a4e34636f72653463686172376d6574686f6473386c656e5f75746638313768343935363635353564666635366333654500656e636f64655f757466385f726177006172697468005f5a4e34345f244c54247538247532302461732475323024636f72652e2e6f70732e2e61726974682e2e52656d244754243372656d313768653539336133626230353330333763654500616c6c6f6300747261697473005f5a4e34636f726535736c6963653469746572313349746572244c54245424475424336e65773137683436326338393130346236666239373745005f5a4e34636f7265336e756d32335f244c5424696d706c24753230247573697a652447542431327772617070696e675f6d756c3137683933396664623563663661656266303945006e6577006d656d6368720077726170005f5a4e34636f726533666d74386275696c6465727331304465627567496e6e657235656e7472793137686361303935346134373764373230616545005f5a4e34636f726533666d74386275696c6465727331304465627567496e6e657235656e74727932385f24753762242475376224636c6f73757265247537642424753764243137686336663430636230393339663733626645005f5a4e34636f726533666d74336e756d313247656e65726963526164697837666d745f696e743137683330323730653937613764383866626145007061640070616e6963005f5a4e34636f726533666d74336e756d35335f244c5424696d706c2475323024636f72652e2e666d742e2e4c6f7765724865782475323024666f7224753230246936342447542433666d74313768663235653065383534373535336437314500696d7000616c7465726e617465006d6170005f5a4e3130325f244c5424636f72652e2e697465722e2e61646170746572732e2e6d61702e2e4d6170244c5424492443244624475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722447542434666f6c643137683439653563633739303661396231626645007772697465007b696d706c23377d006d696e5f62793c7573697a652c20666e28267573697a652c20267573697a6529202d3e20636f72653a3a636d703a3a4f72646572696e673e006765743c267374722c207573697a653e005f5a4e34636f726535736c69636535696e64657837345f244c5424696d706c2475323024636f72652e2e6f70732e2e696e6465782e2e496e646578244c542449244754242475323024666f72247532302424753562245424753564242447542435696e64657831376835623336343435386238326632343635450053706c6974496e7465726e616c006e6578743c636861723e0057726974650077726974655f636861723c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e007b696d706c2332367d005f5a4e34636f72653970616e69636b696e67313870616e69635f6e6f756e77696e645f666d743137683133386130386530383963323036303445005f5a4e34325f244c54242452462454247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d74313768633230363132656137383639386165344500666d74007b696d706c23307d004f7074696f6e007b696d706c23387d005f5a4e34636f726533707472376d75745f70747233315f244c5424696d706c2475323024244250246d757424753230245424475424336164643137686433383935323761353331303836366545006765745f756e636865636b65643c267374723e005f5a4e34636f726533666d7439466f726d6174746572313264656275675f73747275637431376838333134343030643138313466376534450070616e69635f737472005f5a4e34636f726533666d74386275696c64657273313564656275675f7475706c655f6e65773137683134383664383033383865636636373745005553495a455f4d41524b455200736c696365005f5a4e34636f7265336d656d377265706c6163653137683665313530623565366261663964346545007061645f696e74656772616c006765743c75383e005f5a4e34636f726535736c6963653469746572313349746572244c54245424475424336e65773137686231373834333338323430613463363745007b696d706c2331397d006e6578745f6d61746368005f5a4e34636f726536726573756c743139526573756c74244c542454244324452447542438616e645f7468656e3137686639613762303833656534636237383245005f5a4e37335f244c5424636f72652e2e666d742e2e6e756d2e2e5570706572486578247532302461732475323024636f72652e2e666d742e2e6e756d2e2e47656e657269635261646978244754243564696769743137683933663339316566393536306361643245005f5a4e34636f72653370747231303264726f705f696e5f706c616365244c542424524624636f72652e2e697465722e2e61646170746572732e2e636f706965642e2e436f70696564244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c542475382447542424475424244754243137683465633534623435323134663763393045005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683334323336653433336537396333623345006c74006368617273005f5a4e34636f72653373747232315f244c5424696d706c247532302473747224475424336765743137686361316261643162613538333362626645006765743c636f72653a3a6f70733a3a72616e67653a3a52616e6765546f3c7573697a653e3e00706f73745f696e635f73746172743c7573697a653e005f5a4e37355f244c54247573697a65247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c54242475356224542475356424244754242447542431336765745f756e636865636b65643137686630663432666234656339376261626145006164643c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e006d6574686f6473005f5a4e34636f726533666d74386275696c64657273313050616441646170746572347772617032385f24753762242475376224636c6f737572652475376424247537642431376862353032353031383864353564626337450063617061636974795f6f766572666c6f7700666d745f753634005f5a4e36385f244c5424636f72652e2e666d742e2e6275696c646572732e2e50616441646170746572247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f7374723137686539366438303337316562386433343445005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243361646431376836343831303738333031643161616237450049746572005f5a4e34636f72653373747232315f244c5424696d706c2475323024737472244754243563686172733137683635643537336338666664393434333645005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f723130616476616e63655f62793137683837343136383366376333383664636245006e6578745f636f64655f706f696e743c636f72653a3a736c6963653a3a697465723a3a497465723c75383e3e005f5a4e39335f244c5424636f72652e2e736c6963652e2e697465722e2e4368756e6b73244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137686264343939663734373230663065386245004f7264006164643c267374723e007b696d706c23367d00616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23357d3a3a656e7472793a3a7b636c6f737572655f656e7623307d3e004465627567536574005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f666d743137683565373464633863623261616161323645007b696d706c23327d005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542434697465723137686331616261316236653465646465623545005f5a4e34636f726533666d7439466f726d6174746572336e65773137686165623034366666366431666231663445005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243361646431376838353436653232346135313966363633450064656275675f7374727563745f6e657700746f5f7538005f5a4e34636f726533636d7035696d706c7336395f244c5424696d706c2475323024636f72652e2e636d702e2e5061727469616c4571244c54242452462442244754242475323024666f7224753230242452462441244754243265713137683436393566636435376362636161326145005f5a4e34636f726533666d743577726974653137683537653362636463656237646630393145006578706563745f6661696c6564006c656e5f6d69736d617463685f6661696c006f707300696e7472696e736963730073756d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e005f5a4e34636f7265336d656d377265706c61636531376838363534306363336630326138396663450069735f6e6f6e653c7573697a653e00697465723c5b7573697a653b20345d3e00696e746f5f697465723c5b7573697a653b20345d3e005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683366313636623661373436326234373945005f5a4e34636f726533666d7432727438417267756d656e7433666d74313768363232636537653835383430326338654500666d745f696e743c636f72653a3a666d743a3a6e756d3a3a4c6f7765724865782c207536343e00657175616c3c75382c2075383e005f5a4e34636f726535736c696365366d656d63687231326d656d6368725f6e616976653137686363623962373463393862393633336245006d656d6368725f6e6169766500616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23347d3a3a66696e6973683a3a7b636c6f737572655f656e7623307d3e005f5f616c6c6f635f6572726f725f68616e646c657200636f6e73745f707472005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f723373756d313768616537613566613764646461346162384500757466385f69735f636f6e745f62797465006e6578743c636f72653a3a666d743a3a72743a3a417267756d656e743e005f5a4e34636f726533666d74386275696c64657273313664656275675f7374727563745f6e65773137686135363836656238343531653037323245005f5a4e34636f72653970616e69636b696e67313370616e69635f646973706c6179313768663965353336303933393038663832624500656e64735f776974683c636861723e0065713c75382c2075383e007b696d706c23347d005f5a4e34636f726533737472313176616c69646174696f6e733137757466385f69735f636f6e745f6279746531376861396331376363326537313134623836450073706c69745f61745f756e636865636b65643c75383e0073706c69745f61743c75383e005f5a4e34636f72653373747235636f756e74313873756d5f62797465735f696e5f7573697a653137683733663965326535343130353136333245006e6578743c636f72653a3a666d743a3a72743a3a506c616365686f6c6465723e00417267756d656e74005f5a4e37355f244c54247573697a65247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c54242475356224542475356424244754242447542431336765745f756e636865636b6564313768656630633435353430343632353962624500636f6e7461696e735f7a65726f5f62797465005f5a4e37395f244c5424636f72652e2e726573756c742e2e526573756c74244c5424542443244524475424247532302461732475323024636f72652e2e6f70732e2e7472795f74726169742e2e54727924475424366272616e63683137683034646133323232663535363066313845005f5a4e34636f7265366f7074696f6e31336578706563745f6661696c65643137686332333330616533386638616564396545005f5a4e34636f726533707472376d75745f70747233315f244c5424696d706c2475323024244250246d7574247532302454244754243361646431376837336363316163653933303039363536450073756d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e2c207573697a653e005f5a4e35365f244c54247573697a65247532302461732475323024636f72652e2e697465722e2e7472616974732e2e616363756d2e2e53756d244754243373756d32385f24753762242475376224636c6f73757265247537642424753764243137683665653564323561643365666465373945007369676e5f61776172655f7a65726f5f70616400726561643c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e006e6578743c7573697a653e00756e777261705f6f723c267374723e005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243136616c69676e5f746f5f6f6666736574733137683265333033653231353164623038353745005f5a4e34636f726535736c69636532395f244c5424696d706c2475323024247535622454247535642424475424336765743137683037666466393631613031323632356145006e65773c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e007b696d706c2334347d0070616e69635f6e6f756e77696e645f666d740077726974655f7374723c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e577269746524475424313077726974655f636861723137683239666437616639333939643762333645005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243135636f70795f66726f6d5f736c69636531376c656e5f6d69736d617463685f6661696c3137686531663934356265353831313135613845006c6962726172792f616c6c6f632f7372632f6c69622e72732f402f616c6c6f632e643733613839653266303538366464312d6367752e30004974657261746f7200636f756e745f6368617273005f5a4e34636f72653469746572386164617074657273336d6170386d61705f666f6c6432385f24753762242475376224636c6f73757265247537642424753764243137686265643362346664336632356561633645005f5a4e34636f7265366f7074696f6e31354f7074696f6e244c542454244754243769735f6e6f6e653137683036303537623832613939663564313445005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542438616c69676e5f746f3137686361663565313535373365303734303345007b696d706c2331317d005f5a4e34636f726533636d70366d696e5f62793137683961363365346463336265666132393045005f5a4e34636f7265336d656d31326d617962655f756e696e697432304d61796265556e696e6974244c54245424475424357772697465313768643262633963366561386361383161624500656e636f64655f75746638005f5a4e34636f726533666d743557726974653977726974655f666d743137683364623431343565346436363932376245006669656c64007b696d706c2334307d005f5a4e36305f244c5424636f72652e2e63656c6c2e2e426f72726f774572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137686163386261333334363731373261333845005f5a4e34636f726533666d74336e756d35325f244c5424696d706c2475323024636f72652e2e666d742e2e4c6f7765724865782475323024666f72247532302469382447542433666d743137683039663834613031663936303437366145006e6578743c75383e00746f5f7573697a65006d656d005f5a4e34636f7265337074723577726974653137683934303032343231393363646338316545005f5a4e38395f244c5424636f72652e2e6f70732e2e72616e67652e2e52616e6765244c54245424475424247532302461732475323024636f72652e2e697465722e2e72616e67652e2e52616e67654974657261746f72496d706c2447542439737065635f6e65787431376834303038636235396134653064623339450061735f7573697a65006164643c636f72653a3a666d743a3a72743a3a417267756d656e743e00696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e005f5a4e34636f7265336e756d32335f244c5424696d706c24753230247573697a652447542431327772617070696e675f73756231376838643635306338643866353735643162450069735f70726574747900616461707465727300726561643c636861723e007b696d706c23337d00636861725f696e646963657300616c69676e5f746f3c75382c207573697a653e007772617070696e675f6d756c0077726974653c75383e005f5a4e35305f244c5424753634247532302461732475323024636f72652e2e666d742e2e6e756d2e2e446973706c6179496e742447542435746f5f75383137683636316463333963356464386666653545007061747465726e0069735f7375666669785f6f66005f5a4e34636f726535736c696365366d656d63687231346d656d6368725f616c69676e6564313768643864383232303663636532343531614500526573756c740050616441646170746572005f5a4e34636f726533666d7439466f726d6174746572337061643137683433336537613934646232626438653245005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f7374723137683865303931326361326264646233386345005f5a4e34636f726533666d7432727431325553495a455f4d41524b455232385f24753762242475376224636c6f7375726524753764242475376424313768643137376134333532613130653633314500466e4f6e6365006e756d005f5a4e38315f244c5424636f72652e2e7374722e2e697465722e2e4368617273247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722447542435636f756e743137686638633866336432633063356164333545005f5a4e34636f726533666d7439466f726d617474657231397369676e5f61776172655f7a65726f5f7061643137683136323439616566366630343733333545006e65773c75383e007b696d706c23357d005f5a4e34636f726533636d70334f7264336d696e31376861623865636338303366663033636364450072756e005f5a4e34636f726533666d74386275696c64657273313044656275675475706c653969735f7072657474793137683131646663373739346165376162303045005f5a4e34636f726533666d7439466f726d617474657231327061645f696e74656772616c313277726974655f70726566697831376838346635386564303837613362643933450066756e6374696f6e00466f726d61747465720066696c746572006d61705f666f6c64005f5a4e38315f244c5424636f72652e2e7374722e2e697465722e2e4368617273247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683064323235303663643135633337363345007b696d706c2337307d005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683634663237353939353136663335636545005f5a4e35355f244c542424524624737472247532302461732475323024636f72652e2e7374722e2e7061747465726e2e2e5061747465726e24475424313269735f7375666669785f6f663137686536396533336230613062663235373545007772617070696e675f7375620077726974655f666d743c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e005f5a4e35616c6c6f63377261775f766563313763617061636974795f6f766572666c6f7731376837363964333737343539393364316265450063616c6c5f6f6e63653c636f72653a3a666d743a3a72743a3a5553495a455f4d41524b45523a3a7b636c6f737572655f656e7623307d2c2028267573697a652c20266d757420636f72653a3a666d743a3a466f726d6174746572293e0062000000020000000000740000003400000063617061636974795f6f766572666c6f77002f0000007261775f76656300590000005f5f72646c5f6f6f6d004f000000616c6c6f6300540000005f5f616c6c6f635f6572726f725f68616e646c65720000000000f31b0000020074000000282600006a01000077726974653c636861723e00e22100006d617962655f756e696e697400bf2400006272616e63683c28292c20636f72653a3a666d743a3a4572726f723e00e90000006d75745f70747200c0220000696e736572743c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e00070400007b696d706c2334317d00ed1b0000636f70795f6e6f6e6f7665726c617070696e673c75383e005d060000466f726d617474657200ab2300007b696d706c2331377d00cc1f0000737065635f6e6578743c7573697a653e00701c0000706f73745f696e635f73746172743c7573697a653e00a71b0000617269746800d8180000446562756753657400091b00007b696d706c2332357d008d240000526573756c7400e72000006e6578745f636f64655f706f696e743c636f72653a3a736c6963653a3a697465723a3a497465723c75383e3e0034000000726561645f766f6c6174696c653c7573697a653e00151d0000697465723c5b7573697a653b20345d3e00d52100007265706c6163653c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e008d1f00007b636c6f7375726523307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e00e11c000073706c69745f61745f756e636865636b65643c75383e00c82100007265706c6163653c636861723e00a622000069735f6e6f6e653c7573697a653e002f1d00006765743c267374722c207573697a653e000d2500007b696d706c2332367d004321000069735f636861725f626f756e64617279006e240000726573756c7400581b000066756e6374696f6e00831f0000636f756e7400960600007061645f696e74656772616c00fb1c0000616c69676e5f746f5f6f6666736574733c75382c207573697a653e00751d00006c656e5f6d69736d617463685f6661696c00da0000006164643c75383e00581c00006e65773c75383e00fa030000646967697400211b0000666d743c28293e005523000070616e69636b696e6700b3220000756e777261705f6f723c267374723e0061200000636f6e7461696e735f6e6f6e5f636f6e74696e756174696f6e5f6279746500cd000000616c69676e5f6f66667365743c75383e00a71c00006e65773c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e000c2400007b696d706c2331397d00462300007772617070696e675f737562006f060000616c7465726e61746500322200006c74005a1f00006d61705f666f6c64006d20000073756d5f62797465735f696e5f7573697a6500ae010000417267756d656e7400e72100004d61796265556e696e6974009a050000666d7400b11b000072656d00ce2200006578706563745f6661696c656400f1020000666d745f696e743c636f72653a3a666d743a3a6e756d3a3a4c6f7765724865782c2075383e00bb1e0000636f6e7461696e735f7a65726f5f62797465004f13000072756e00c22000007b696d706c2334347d00882100007b696d706c2332387d003313000077726974655f707265666978005d1b0000466e4f6e636500da1d00006765743c267374723e005b000000636f6e73745f70747200b32100006e6578745f6d6174636800631d00006765743c75382c20636f72653a3a6f70733a3a72616e67653a3a52616e67653c7573697a653e3e00e5020000666d745f696e743c636f72653a3a666d743a3a6e756d3a3a55707065724865782c2075383e001322000077726974653c75383e00340100006164643c7573697a653e00471c00004974657200dd14000064656275675f7374727563745f6e6577001c1b00007b696d706c2335337d00b30000006164643c636f72653a3a666d743a3a72743a3a417267756d656e743e0009200000737472007323000070616e69635f646973706c61793c267374723e00ba1c0000697465723c75383e00701d0000636f70795f66726f6d5f736c69636500431f00006d617000832100007061747465726e00d9020000666d745f696e743c636f72653a3a666d743a3a6e756d3a3a4c6f7765724865782c207536343e005617000066696e69736800f50300007b696d706c2332397d00ac240000616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23347d3a3a66696e6973683a3a7b636c6f737572655f656e7623307d3e0073240000756e777261705f6661696c6564000a1c00006e6578743c75383e00af20000053706c6974496e7465726e616c003d200000646f5f636f756e745f6368617273003a1c00006e6578743c636f72653a3a666d743a3a72743a3a417267756d656e743e00fb1b0000736c696365006a17000044656275675475706c6500881f0000746f5f7573697a65004c1c0000706f73745f696e635f73746172743c75383e007a2000006974657200291f000073756d002d2200007b696d706c2335347d007d1c00007b696d706c2337307d00ce1d00006765745f756e636865636b65643c636f72653a3a666d743a3a72743a3a417267756d656e743e009f240000616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23357d3a3a656e7472793a3a7b636c6f737572655f656e7623307d3e00551a00007b696d706c23307d002b200000636861725f636f756e745f67656e6572616c5f6361736500a021000069735f7375666669785f6f66004d1f0000666f6c643c7573697a652c20636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c207573697a652c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e0025120000777261705f6275663c636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23317d3a3a777261703a3a7b636c6f737572655f656e7623307d3e00da1a000077726974655f666d743c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e00e3010000666d745f753634002a000000636f726500081d000061735f6368756e6b733c7573697a652c20343e000813000064656275675f7475706c655f6669656c64315f66696e697368009c0100005553495a455f4d41524b4552003e1f00006164617074657273002c2300007772617070696e675f6d756c002e1f00007b636c6f7375726523307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e004f2100006765743c636f72653a3a6f70733a3a72616e67653a3a52616e6765546f3c7573697a653e3e00a60000006164643c5b7573697a653b20345d3e00771f0000636f756e743c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e00951c0000696e746f5f697465723c5b7573697a653b20345d3e00dd1e0000666f6c643c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a6d61703a3a6d61705f666f6c643a3a7b636c6f737572655f656e7623307d3c2675382c207573697a652c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e3e00871800007b696d706c23317d008b23000070616e69635f6e6f756e77696e645f666d7400ed25000063686172006d1f000066696c746572009d1f0000656e756d657261746500971e00006d656d6368725f6e61697665008906000070616464696e67002e0300007b696d706c2336347d00181f00007b696d706c2334387d008c1800007772617000ca19000064656275675f7475706c655f6e657700e91400007b696d706c23327d00b301000061735f7573697a65001d1f000073756d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e0028220000696d706c7300ac1b00007b696d706c233232357d00131f0000616363756d00d81900005772697465005a23000070616e6963002e1c00006e6578743c636f72653a3a666d743a3a72743a3a506c616365686f6c6465723e0029210000636861727300531b00006f707300f22500006d6574686f647300781e000065713c75382c2075383e00c72000006e6578743c636861723e00950500007b696d706c2336357d005c210000656e64735f776974683c636861723e00c32100006d656d009b2100007b696d706c23337d007f23000070616e69635f737472007c1700006669656c64006e2200004f72640097010000727400de010000696d7000a71f00006e6578743c636f72653a3a736c6963653a3a697465723a3a497465723c636f72653a3a666d743a3a72743a3a506c616365686f6c6465723e3e00221c00006e6578743c7573697a653e00a21c0000497465724d75740069130000777269746500491d0000656e64735f776974683c75383e00b118000069735f70726574747900161c00006e6578743c5b7573697a653b20345d3e009f1800004465627567496e6e657200dd180000656e74727900f71e0000616476616e63655f62793c636f72653a3a7374723a3a697465723a3a43686172496e64696365733e00d402000047656e657269635261646978006a21000074726169747300fd020000666d745f696e743c636f72653a3a666d743a3a6e756d3a3a55707065724865782c207536343e005a1a000077726974655f7374723c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e00a22000006e65787400ea1e000073756d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e2c207573697a653e003e1700007b696d706c23347d00ee14000077726974655f73747200f72500006c656e5f75746638005222000065713c5b75385d2c205b75385d3e005d010000726561643c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e00ee1c000073706c69745f61743c75383e00b42000006e6578745f696e636c75736976653c636861723e001c0300007b696d706c2331317d0050010000726561643c636861723e007f090000706164005f1f00007b636c6f7375726523307d3c2675382c207573697a652c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e00731a000077726974655f636861723c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e00f3200000757466385f66697273745f6279746500bf1800007b696d706c23357d00b31f00006e6578743c636f72653a3a736c6963653a3a697465723a3a497465723c636f72653a3a666d743a3a72743a3a417267756d656e743e3e00612200006d696e5f62793c7573697a652c20666e28267573697a652c20267573697a6529202d3e20636f72653a3a636d703a3a4f72646572696e673e00ff1100006e657700152300006e756d007701000077726974653c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e00b81d0000696e64657800942200004f7074696f6e009922000069735f736f6d653c7573697a653e00d81400006275696c646572730036210000636861725f696e646963657300a623000063656c6c00c00000006164643c267374723e00c71c00006765743c75382c207573697a653e00f31d00007b696d706c23367d00411e00006765743c75383e005b1700007b636c6f7375726523307d00db200000757466385f69735f636f6e745f6279746500d81e00004974657261746f7200621b000063616c6c5f6f6e63653c636f72653a3a666d743a3a72743a3a5553495a455f4d41524b45523a3a7b636c6f737572655f656e7623307d2c2028267573697a652c20266d757420636f72653a3a666d743a3a466f726d6174746572293e00a31e00006d656d6368725f616c69676e656400d41c0000616c69676e5f746f3c75382c207573697a653e00221d00006765745f756e636865636b65643c636f72653a3a666d743a3a72743a3a417267756d656e742c207573697a653e00410100006164643c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e00aa1d0000697465725f6d75743c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e008f2200006f7074696f6e0004260000656e636f64655f757466385f72617700d620000076616c69646174696f6e7300501e0000636d70007421000067657400e61d00006765745f756e636865636b65643c267374723e00291300007b696d706c23377d00051c00007b696d706c233138317d00d31e00006974657261746f72001812000064656275675f737472756374002f1e0000696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e2c20636f72653a3a6f70733a3a72616e67653a3a52616e676546726f6d3c7573697a653e3e00041f00006e74683c636f72653a3a7374723a3a697465723a3a43686172496e64696365733e0016260000656e636f64655f75746638007518000050616441646170746572008b1e00006d656d636872006f2100007b696d706c23387d00c11b0000696e7472696e7369637300ff240000696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e2c20636f72653a3a6f70733a3a72616e67653a3a52616e676546726f6d3c7573697a653e2c203132383e00c21f000072616e676500d32400007b696d706c2331357d007c0600007369676e5f61776172655f7a65726f5f70616400620600007369676e5f706c7573002f000000707472004100000064726f705f696e5f706c6163653c26636f72653a3a697465723a3a61646170746572733a3a636f706965643a3a436f706965643c636f72653a3a736c6963653a3a697465723a3a497465723c75383e3e3e001f200000636f756e745f636861727300641c00006e65773c5b7573697a653b20345d3e0016130000506f737450616464696e670017210000757466385f6163635f636f6e745f6279746500f81d0000696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e00402200007b696d706c23397d005c130000676574636f756e740092240000616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23347d3a3a6669656c643a3a7b636c6f737572655f656e7623307d3e00812200006d696e3c7573697a653e0021030000746f5f753800ce0400007b696d706c2334307d005a1e0000657175616c3c75382c2075383e00ce240000617272617900000000000e00000002000000000074000000000000000e0000000200740000002826000000000000412a000000726973637600012000000004100572763634693270305f6d3270305f613270305f633270300084000000040040000000010101fb0e0d0001010101000000010000016c6962726172792f616c6c6f632f73726300007261775f7665632e727300010000616c6c6f632e72730001000000000902326e010000000000038a040105050a030109020001090c000001010402000902406e010000000000038d0301050d0a030b09020001090c00000101781e000004005e030000010101fb0e0d0001010101000000010000016c6962726172792f636f72652f7372632f6f7073006c6962726172792f636f72652f7372632f707472006c6962726172792f636f72652f7372632f666d74006c6962726172792f636f72652f737263006c6962726172792f636f72652f7372632f736c6963652f69746572006c6962726172792f636f72652f7372632f697465722f747261697473006c6962726172792f636f72652f7372632f737472006c6962726172792f636f72652f7372632f69746572006c6962726172792f636f72652f7372632f697465722f6164617074657273006c6962726172792f636f72652f7372632f6d656d006c6962726172792f636f72652f7372632f6d6163726f73006c6962726172792f636f72652f7372632f736c696365006c6962726172792f636f72652f7372632f6e756d006c6962726172792f636f72652f7372632f6172726179006c6962726172792f636f72652f7372632f63686172000066756e6374696f6e2e7273000100006d6f642e72730002000072742e7273000300006e756d2e727300030000636f6e73745f7074722e727300020000696e7472696e736963732e7273000400006d75745f7074722e7273000200006d6f642e7273000300006d6163726f732e7273000500006974657261746f722e72730006000076616c69646174696f6e732e727300070000616363756d2e727300060000636d702e72730004000072616e67652e7273000800006d61702e72730009000066696c7465722e727300090000636f756e742e727300070000697465722e7273000700006d6f642e7273000a00006f7074696f6e2e7273000400006d6f642e7273000b00006d6f642e727300070000696e6465782e7273000c00007472616974732e7273000700006d6f642e7273000c000075696e745f6d6163726f732e7273000d0000697465722e7273000c000070616e69636b696e672e727300040000656e756d65726174652e72730009000063656c6c2e7273000400006275696c646572732e727300030000726573756c742e7273000400006d617962655f756e696e69742e7273000a00006d6f642e7273000e0000636d702e7273000c00007061747465726e2e7273000700006d656d6368722e7273000c00006d6574686f64732e7273000f000061726974682e727300010000000009022ab301000000000003f90101040205090a03860a090000010403050503d3750902000109020000010104020009022eb301000000000003ea030105010a030009000001090200000101040400090230b301000000000003d2010105170a03130906000106039a7e0918000103e60109040001039a7e0924000105150603e80109020001051e0302090e00010405050d03b505091a00010406050903d20d090200010404051e03fa6c0904000104060509038613090400010405050d03ae72090800010406050903d20d090200010404051503fb6c09080001040605090385130902000106030009040001040405170603f56c0908000106039a7e0906000105140603f901090400010515030209040001051e037f091c000105150302090400010405050d03a305090200010406050903d20d090200010407050d039c73090c00010406050903e40c0902000106038f6b090a000104040514060381020902000105150301090400010407050d038b06090800010404051503f67909020001051e0302090a000105150301090200010405050d039905090400010406050903d20d090200010407050d039c73090c00010406050903e40c0902000106038f6b090800010407050d06038d08090400010404053e03827a09060001050d030209020001050a030109140001060b030009020001090400000101040800090272b401000000000003dd090105090a03e003091e0001051303a77c090c000106039b76090c000105090603f70d09040001051303ee7b0904000105190305090200010603967609020001050f0603fb0909020001050906030009020001038576090400010409051806038601090200010603fa7e09040001040a05150603b113090400010407050d03dc7409040001040b0505038c78090200010409051803ed0009080001040c051c03af7f090200010409051803d100090200010408050d03e50809020001050f031009020001050906030009020001052306030909020001051a06030009040001050906038d0409040001051a03f97b09020001051b03e90009020001053103a47f09060001051503dc000904000106038d7509060001050606039d0a09200001060b0300091c0001050003e3750904000104020509060394090926000106030009060001040805110603f900090400010402050903cd00090a000106030009040001040805110603b37f090400010603f3750914000105090603800b09020001040d05340353090600010408050d032e090400010603ff740910000105150603f30a090200010530030a0904000105230603000904000105300300090200010383750906000105090603800b090c0001040d0534035309040001040e050c039a7a090200010408050d039406090200010603ff74090c000105240603970a090a00010511030109040001030109140001050903fb7e090e0001040d053403bf01090800010408050d03c27e09080001051103fa00091000010603f175091000010603910a090200010301090400010603ee7509080001040d05340603d30a09020001090600000101040800090256b601000000000003f2090105140a0301091c0001051103010904000105140302090e0001052c060300090200010b03000912000103897609040001050a0603f80909020001060b0300090a00010904000001010408000902acb601000000000003bb0a01041405120a039b7a090200010408050c03e7050916000104150509039a78090200010408050c03e607090800010518030509040001051d060300090400010405050d0603dc7c09040001040a050903b87b09040001040b05000603a97d09120001041205260603910109040001051106030009020001040a05100603c70109040001040d053403fb0709040001040e050c039a7a090200010409051803997c09020001040b050d03a07f0904000105080301090800010516030a090400010505035b0904000105110306090400010508032109040001051a0305090400010505035a090400010511060300090200010505030009040001050c06032909040001051e030509040001051203010904000105050351090400010511060300090200010505030009040001050d06032f090400010412050903cb00090200010603f47e090400010409051806038601091e0001040b050d03a07f090400010508030109040001060359090400010603330908000106034d09040001050c06033b09040001050006034509040001051a060338090400010511035a0904000106030009040001051e06032e09040001051203010904000105050351090400010511060300090600010505030009040001050d06032f090200010412050903cb00090600010416050c03cc000904000105090304090200010417050c037d0904000104160513030f0904000104180509032c090800010603ec7d0904000104140603bc0709020001041803d87a090400010603ec7d0904000104140603bc07090200010603c4780902000104080603d40a0904000105120304090400010411050803c37509080001060365090400010409051806038601090200010603fa7e09040001040a05150603b113090400010407050d03dc7409040001040b0505038c78090200010409051803ed0009080001040c051c03af7f090200010409051803d100090200010402051f03bb0c0904000104190545036509060001051603800e090800010409051803e065090600010603fa7e09040001040a05150603b113090200010407050d03dc7409040001040b0505038c78090200010409051803ed0009080001040c051c03af7f090200010409051803d100090200010603fa7e090200010386010902000103fa7e09020001040a05150603b113090600010407050d03dc7409040001040b0505038c78090200010409051803ed0009080001040c051c03af7f090200010409051803d100090200010603fa7e09020001041105150603c7000922000105000603b97f09060001051b0603fe00090e00010534060300090400010533030009020001051b030009040001041a050d0603e7080902000104110505039a77090400010509035b09020001050c030609020001041b03e80a090200010603b874090200010419053806039908091200010405050d03867f090400010409051803e779090600010603fa7e09020001041105190603d0000904000105120301090200010507032309020001050606030009040001051203000902000106035d09020001050503230902000105110360090400010507032009020001050606030009040001051206035d090200010323090200010505060300090200010507030009040001050603000904000105120300090200010505030009020001051206035d0902000105050323090200010511036009020001050703200904000105060603000904000105120300090200010505030009020001040905180603120904000104110511034e09040001040905180332090200010603000906000103fa7e090400010386010904000103fa7e09040001038601090600010411051206035d090600010407050d03aa07090200010411050703e7780902000105060603000904000105120300090200010505030009020001040905180603120904000104110511035e09020001040905180322090200010603fa7e090400010411051b0603fe00090200010534060300090400010533030009020001051b030009040001041a050d0603e7080902000104110505039a7709040001050d0367090200010408051403f60909020001051b0317090400010535037009060001051503100904000106038d750906000103f30a09260001053006030a0904000105230603000904000105300300090200010383750906000105090603800b090e0001040d0534035309040001040e050c039a7a090200010408050d039406090200010603ff74090c000105280603e30a090a00010515030109040001050903b07e090e0001040d053403bf0109080001040e050c039a7a090400010408050d03a804090400010603eb7609100001040d05340603d30a0902000104080506031609040001060b030009140001090400000101041c00090224ba01000000000003ed000105050a030709020001090c00000101040800090232ba01000000000003b7080105090a03bb7909180001050b03c90609080001050903b77909040001050503c90609080001050e030e090200010409051803bc78090400010603fa7e0904000103860109040001040805150603cb0709220001051406030009020001051506030109020001052d0603000904000105150300090400010510060313090600010505060300090200010511060301090200010505060300090400010511060301090400010533036f09020001050503110904000105150304090200010505030f090600010403050c039978090600010603ed7e090a0001051d0603960109040001051b0603000902000103ea7e09020001040805090603eb080902000105190301090400010505030e090800010403050c039978090600010603ed7e090a0001051d0603960109040001051b0603000902000103ea7e09020001040805090603ec0809020001052d0307090400010405050d03ac7e090200010403050903eb7909040001051a060300090200010509030009020001040805110603cc07090400010409051803b078090200010408051d03b907091000010409051803c778090400010603fa7e0904000103860109080001040805150603bd0709120001051406030009020001051506030109020001052d060300090400010515030009040001040305090603c67809060001051a060300090200010509030009040001040805110603bc07090400010409051803c078090200010408051a03d707090a00010417050c03fc78090400010603a77e090600010408051a0603dd08090200010417050c03fc78090400010408051a038407090400010405050d03c27e090400010408050903bf0109040001052106030009040001050903000908000103a2770906000105020603e20809060001060b030009100001090400000101041e000902b0bb01000000000003ba0501040805090a03ba0609000001091200000101041e000902c2bb01000000000003d50501040805090a039f06090000010912000001010420000902d4bb01000000000003f10c0105050a030109020001090c000001010414000902e2bb010000000000038a0f01041c05050a038b7209020001090c00000101041c000902f0bb01000000000003cf0001050e0a031009020001090c000001010404000902febb010000000000039901010407050d0a03f30609060001040405000603f3770908000106039301090800010421050903d602090200010404051403ea7c090400010603ad7f09080001052306032a0902000103e900090800010603ed7e090400010417050c0603ed03090a00010404050903817d090a0001050e032e09160001060b0300090200010417050d0603d20209040001090e00000101041f0009026ebc010000000000031e010412050c0a03ce040946000104190523039c0d091800010423050d03d26e09040001041f034a090a00010301090400010412050c03c704090e00010424051903b17e090800010417050c0342090a00010425050803cb7d09080001050b030d0906000106034809040001050c0603390902000105090304090c0001050b037b090200010402051f03890d09060001051b03010908000104250508039273090400010603ac7f090e000105100603eb00090600010405050d03b406090400010425051503c679090400010529030409060001041a050d03e508090200010425050503c67609020001051503d2000908000105290304090a0001041a050d03e408090200010425050503c67609020001050903db0009080001050b037209020001050c03580906000105090304090c0001050b037b09020001060348090400010603e1000904000106039f7f09040001050c06033909060001050b037f090c000106034809080001042405200603b403090200010511060300090200010417050c0603ac7f090800010423050d03fb7d090200010424051c03dd02090400010603c87c09040001041f051006032109140001051103010906000106035e090e00010419050906038912090800010603f76d09040001041f050606032a09100001060b0300091a000109040000010104080009022abe01000000000003a20101052b0a0301090c00010426050803f60b09020001050d031f09040001050f0363090800010513032009060001050d06030009040001051206030109080001050d06030009040001050f060361090c00010513032209060001050d06030009040001051206030109080001050d06030009060001051206030109080001050d060300090400010512060303090c0001050d06030009060001051206030109080001050d06030009060001051206030109080001050d06030009060001051206030109080001050d06030009040001040805090603dc73090a000105060301090a0001060b0300090200010904000001010408000902debe01000000000003be010105090a0301090200010506030109300001060b030009020001090400000101040800090216bf01000000000003c5010105090a030109000001090a00000101040800090220bf01000000000003c9010105090a030109020001052b0359090c00010426050803f60b09020001050d031f09040001050f0363090800010513032009060001050d06030009040001051206030109080001050d06030009040001050f060361090c00010513032209060001050d06030009040001051206030109080001050d06030009060001051206030109080001050d060300090400010512060303090c0001050d06030009060001051206030109080001050d06030009060001051206030109080001050d06030009060001051206030109080001050d06030009040001040805090603dc73090a000105060328090a0001060b0300090200010904000001010408000902d6bf01000000000003cd010105090a0301090200010371091e00010506031009140001060b030009020001090400000101041f00090210c001000000000003b3020105170a0301091200010420050903f10709040001041f03a078090200010603ba7d0908000105100603b602090400010408050903c10b09040001041f050006038972090400010408050903f70d09040001041f05100603bf740904000105000603ca7d09020001051e0603c002090400010603c07d0904000105140603b702090a00010408050903be0909040001041f051503c376091600010603c87d09020001040805090603f50b090e0001041f051e03cb76090a00010408050903b50909020001042003a70309040001041f051103a673090200010408051403e406090c00010603da7609040001041f05210603bb02090200010408051703e806090400010414050903f002090800010408051303947d090a0001051403010904000103010904000105180301090800010509037709080001041f0511039c79091400010408050903e40609040001041f0511039c79090a00010408050903b80909080001041f050006038b740912000105090603b502090200010311090400010506030209060001060b030009100001090400000101041f00090230c101000000000003d3030105170a03a87f091200010420050903aa0709080001041f03d67809020001031209040001050603c90009040001060b03000910000103a97c0904000105100603fd02090400010408050903fa0a09040001041f050006038972090400010408050903f70d09040001041f051006038675090400010514030a090200010408050903ee0809020001041f051503937709180001051103020902000105140374090a00010408050903f70809020001041f0515038a77091800010408051403a706090200010603da7609040001041f052106038203090200010408051703a106090400010414050903f002090800010408051303947d090a0001051403010904000103010904000105180301090800010509037709080001041f051103e379091e00010408050903f10809080001091600000101040800090230c201000000000003e40f0105090a03907c090c0001041f050503a376090c00010408050903cf0d090c0001041f050c03fd72090e0001050006039c7d09020001050c03e40209040001039c7d09020001042005090603a60a09020001041f051403c07809020001050006039a7d090a0001051403e60209020001040805090603910b09080001041f051403ef740906000104080509038f0909020001041f051503f2760914000104080509038e0909020001041f03f776091600010408050603fd0c09040001060b0300090a00010904000001010419000902c8c2010000000000038a1a01050d0a030109020001090c000001010404000902d6c2010000000000039901010407050d0a03f30609060001040405000603f3770908000106039401090c00010421050903d502090200010404051403ea7c090400010427052d03ef03090800010404052303d27c090800010603ec7e090400010417050c0603ed03090a00010404050903817d090a0001050e032e09160001060b0300090200010417050d0603d20209040001090e00000101040400090248c3010000000000039901010407050d0a03f30609060001040405000603f3770908000106039301090c00010421050903d602090200010404051403ea7c090400010427052d03ef03090800010404052303d17c090800010603ed7e090400010417050c0603ed03090a00010404050903817d090a0001050e032e09160001060b0300090200010417050d0603d20209040001090e000001010408000902bac301000000000003cf110105090a03ec01090000010916000001010422000902d0c301000000000003820101040805090a03f20a090a00010422051e038f75090200010408050903f10a09020001041f050503a376091000010408050903cf0d090c0001041f050c03fd7209140001050006039c7d09020001050c03e40209040001039c7d09020001042005090603a60a09020001041f051403c07809020001050006039a7d090a0001051403e60209020001040805090603910b09080001041f051403ef740906000104080509038f0909020001041f051503f2760914000104080509038e0909020001041f03f776091600010422050f03977e09040001060b030009080001090400000101040400090272c4010000000000039901010407050d0a03f30609060001040405000603f3770908000106039401090800010421050903d502090200010404051403ea7c090400010603ad7f09080001052306032a0902000103ea00090800010603ec7e090400010417050c0603ed03090a00010404050903817d090a0001050e032e09160001060b0300090200010417050d0603d20209040001090e00000101004743433a2028292031322e322e30004c696e6b65723a204c4c442031362e302e320000000000000000000000000000000000000000000000000000000000000000010000000400f1ff00000000000000000000000000000000220000000000050038c902000000000000000000000000002b000000020004008a36010000000000640000000000000000000000000004008a36010000000000000000000000000000000000000004008c360100000000000000000000000000000000000000040094360100000000000000000000000000fc00000000000400a0360100000000000000000000000000080100000200040086c801000000000056000000000000006701000002000400106e01000000000008000000000000000000000000000400ee3601000000000000000000000000007601000002000400ee3601000000000010000000000000000000000000000400ee3601000000000000000000000000000000000000000400fe360100000000000000000000000000c701000002000400fe36010000000000ee000000000000000000000000000400fe36010000000000000000000000000000000000000004000037010000000000000000000000000000000000000004000a3701000000000000000000000000004202000000000400d63701000000000000000000000000004e02000001000100e2090100000000002b00000000000000780200000200040024ba0100000000000e000000000000000000000000000400ec370100000000000000000000000000a502000002000400ec37010000000000d4040000000000000000000000000400ec3701000000000000000000000000000000000000000400ee370100000000000000000000000000000000000000040008380100000000000000000000000000f8020000020004001a47010000000000c600000000000000ce03000002000400043e01000000000030000000000000001f04000002000400343e01000000000030000000000000007404000002000400283d010000000000dc000000000000008f05000000000400563c01000000000000000000000000009b05000001000100690b0100000000003500000000000000c605000000000400643c0100000000000000000000000000d205000001000100410b0100000000002800000000000000fd05000002000400c8c20100000000000e0000000000000063060000000004007a3c01000000000000000000000000006f06000000000400903c01000000000000000000000000007b060000000004009e3c01000000000000000000000000008706000000000400a83c01000000000000000000000000009306000001000100f00a0100000000003000000000000000be06000000000400b63c01000000000000000000000000000000000000000400c03c0100000000000000000000000000ca06000002000400c03c01000000000068000000000000000000000000000400c03c01000000000000000000000000009207000002000400f0bb0100000000000e000000000000000000000000000400283d01000000000000000000000000000000000000000400283d010000000000000000000000000000000000000004002a3d01000000000000000000000000000000000000000400403d01000000000000000000000000000000000000000400043e01000000000000000000000000000000000000000400043e01000000000000000000000000000000000000000400063e01000000000000000000000000000000000000000400083e0100000000000000000000000000cd07000002000400086e0100000000000800000000000000da07000002000400286e0100000000000a000000000000000000000000000400343e01000000000000000000000000000000000000000400343e01000000000000000000000000000000000000000400363e01000000000000000000000000000000000000000400383e01000000000000000000000000000000000000000400643e0100000000000000000000000000f507000002000400643e0100000000007a010000000000000000000000000400643e01000000000000000000000000000000000000000400663e010000000000000000000000000000000000000004007e3e01000000000000000000000000005b08000000000400a23f01000000000000000000000000006708000001000100b90b01000000000033000000000000009208000000000400b03f01000000000000000000000000009f08000001000100ec0b0100000000002700000000000000ca08000000000400be3f0100000000000000000000000000d708000000000400c83f0100000000000000000000000000e408000001000100130c01000000000028000000000000000000000000000400de3f01000000000000000000000000000f09000002000400de3f010000000000aa010000000000000000000000000400de3f01000000000000000000000000000000000000000400e03f01000000000000000000000000000000000000000400fa3f010000000000000000000000000076090000000004005041010000000000000000000000000083090000010001003b0c0100000000003200000000000000ae090000000004005e410100000000000000000000000000bb090000010001006d0c0100000000002800000000000000e60900000000040068410100000000000000000000000000f30900000000040072410100000000000000000000000000000000000000040088410100000000000000000000000000000a0000020004008841010000000000c00100000000000000000000000004008841010000000000000000000000000000000000000004008a4101000000000000000000000000000000000000000400a4410100000000000000000000000000700a000000000400244301000000000000000000000000007d0a000001000100950c0100000000009100000000000000a80a00000000040032430100000000000000000000000000b50a000001000100260d0100000000002a00000000000000000000000000040048430100000000000000000000000000e00a0000020004004843010000000000820100000000000000000000000004004843010000000000000000000000000000000000000004004a4301000000000000000000000000000000000000000400644301000000000000000000000000003e0b000000000400b44401000000000000000000000000000000000000000400ca4401000000000000000000000000004b0b000002000400ca4401000000000050020000000000000000000000000400ca4401000000000000000000000000000000000000000400cc4401000000000000000000000000000000000000000400e644010000000000000000000000000000000000000004001a47010000000000000000000000000000000000000004001a47010000000000000000000000000000000000000004001c4701000000000000000000000000000000000000000400344701000000000000000000000000000000000000000400e04701000000000000000000000000000000000000000400e04701000000000000000000000000000000000000000400e447010000000000000000000000000000000000000004001848010000000000000000000000000000000000000004001848010000000000000000000000000000000000000004001a480100000000000000000000000000990c0000000004001a480100000000000000000000000000a60c00000100060088ca0200000000001000000000000000cf0c0000020004002cae010000000000c204000000000000080d00000200040006b301000000000024000000000000003f0d0000020004004c380200000000001c00000000000000b20d0000020004006838020000000000da00000000000000e80d0000020004007ac60100000000004e00000000000000300e000002000400204a0200000000008601000000000000710e0000020004004aac0100000000008200000000000000b20e000002000400243802000000000028000000000000002b0f000000000400824f0100000000000000000000000000380f0000010001000c050100000000001100000000000000640f000000000400c84f0100000000000000000000000000710f00000200040010aa010000000000c001000000000000a90f00000000040022500100000000000000000000000000b60f00000200040060930100000000007c00000000000000f80f000000000400ee5001000000000000000000000000000510000002000400daa901000000000036000000000000005f100000000004009a5101000000000000000000000000006c10000000000400d851010000000000000000000000000079100000000004000452010000000000000000000000000086100000000004001e5201000000000000000000000000009310000001000100d00401000000000021000000000000009c10000002000400faa30100000000002200000000000000171100000200040088a1010000000000d600000000000000ab110000020004001ca40100000000003a00000000000000e41100000200040052a501000000000042000000000000002312000000000400b25201000000000000000000000000003012000000000400ca5201000000000000000000000000003d12000001000100b0050100000000001c000000000000004712000000000400f0520100000000000000000000000000541200000200040056a4010000000000fc00000000000000dc120000020004008ea30100000000006c000000000000000f1300000200040058a6010000000000640000000000000062130000020004000e5002000000000054020000000000009a1300000200040058720100000000005800000000000000fa13000002000400fc4d0200000000009a000000000000002c140000020004005e7001000000000058000000000000008314000002000400ae6f0100000000005800000000000000df1400000200040006700100000000005800000000000000391500000200040042390200000000002a020000000000006e15000002000400fe6e0100000000005800000000000000cb15000002000400566f01000000000058000000000000002616000002000400b670010000000000580000000000000081160000020004004e6e0100000000005800000000000000dc16000002000400a66e01000000000058000000000000003517000002000400d4a801000000000072000000000000008b170000020004005ccf010000000000ba000000000000000c180000020004000e71010000000000520000000000000065180000020004009e3b02000000000018030000000000009c18000002000400da730100000000004e00000000000000fd180000020004000873010000000000860000000000000049190000020004008e730100000000004c000000000000009519000002000400b0720100000000005800000000000000e01900000200040060710100000000005800000000000000331a00000200040028740100000000009400000000000000941a000002000400d4590200000000007400000000000000c21a000002000400485a0200000000004a3a000000000000f61a000002000400d2450200000000004e04000000000000321b000002000400b8710100000000005200000000000000921b000002000400b63e0200000000008c03000000000000d61b0000020004000a720100000000004e00000000000000291c0000020004006ed1010000000000c000000000000000b51c00000200040062520200000000007207000000000000f41c000002000400424202000000000090030000000000003b1d000002000400964e0200000000007801000000000000701d000002000400bc740100000000009400000000000000d11d000000000400ba6c0100000000000000000000000000de1d000000000400ca6c0100000000000000000000000000eb1d00000100010000020100000000001c00000000000000f11d000000000400d66c0100000000000000000000000000fe1d0000010001005e0a0100000000002b00000000000000291e000000000400de6c0100000000000000000000000000361e00000100010040020100000000002000000000000000601e000002000400d4bb0100000000000e00000000000000931e000000000400f66c0100000000000000000000000000a01e000000000400026d0100000000000000000000000000ad1e000000000400146d0100000000000000000000000000ba1e0000000004001c6d0100000000000000000000000000c71e00000100010020020100000000002000000000000000f11e0000000004002e6d0100000000000000000000000000fe1e000000000400366d01000000000000000000000000000b1f000000000400406d0100000000000000000000000000181f000000000400486d0100000000000000000000000000251f000000000400526d0100000000000000000000000000321f0000000004005a6d01000000000000000000000000003f1f000000000400646d01000000000000000000000000004c1f000001000100200b01000000000021000000000000000000000000000400706d0100000000000000000000000000771f000002000400706d0100000000000a000000000000000000000000000400706d0100000000000000000000000000891f000002000400eeb2010000000000180000000000000000000000000004007a6d0100000000000000000000000000be1f0000020004007a6d010000000000080000000000000000000000000004007a6d0100000000000000000000000000c91f000002000400c299010000000000d4030000000000000000000000000400826d01000000000000000000000000005420000002000400826d01000000000008000000000000000000000000000400826d01000000000000000000000000006120000002000400969d010000000000f20300000000000000000000000004008a6d0100000000000000000000000000ee200000020004008a6d0100000000004e0000000000000000000000000004008a6d010000000000000000000000000000000000000004008c6d01000000000000000000000000000000000000000400966d01000000000000000000000000000000000000000400d86d0100000000000000000000000000fb20000002000400d86d01000000000030000000000000000000000000000400d86d01000000000000000000000000000000000000000400da6d01000000000000000000000000000000000000000400e06d01000000000000000000000000000000000000000400086e01000000000000000000000000000000000000000400086e01000000000000000000000000000000000000000400106e01000000000000000000000000000000000000000400106e01000000000000000000000000000000000000000400186e01000000000000000000000000000d21000002000400186e01000000000008000000000000000000000000000400186e01000000000000000000000000000000000000000400206e01000000000000000000000000001c21000002000400206e01000000000008000000000000000000000000000400206e01000000000000000000000000000000000000000400286e01000000000000000000000000000000000000000400286e01000000000000000000000000003021000002000400406e0100000000000e000000000000000000000000000400326e01000000000000000000000000003a21000002000400326e0100000000000e000000000000000000000000000400326e01000000000000000000000000000000000000000400326e01000000000000000000000000000000000000000400326e01000000000000000000000000000000000000000400346e01000000000000000000000000000000000000000400346e01000000000000000000000000000000000000000400366e01000000000000000000000000000000000000000400406e01000000000000000000000000000000000000000400406e01000000000000000000000000000000000000000400406e01000000000000000000000000000000000000000400406e01000000000000000000000000000000000000000400406e01000000000000000000000000000000000000000400426e01000000000000000000000000000000000000000400426e01000000000000000000000000000000000000000400446e010000000000000000000000000000000000000004004e6e010000000000000000000000000000000000000004004e6e010000000000000000000000000000000000000004004e6e01000000000000000000000000000000000000000400506e01000000000000000000000000000000000000000400546e0100000000000000000000000000732100000200040080cb0100000000006601000000000000ba2100000200040040ce010000000000a2000000000000005722000000000400866e010000000000000000000000000064220000000004008e6e01000000000000000000000000007122000001000100600201000000000020000000000000000000000000000400a66e01000000000000000000000000000000000000000400a66e01000000000000000000000000000000000000000400a86e01000000000000000000000000000000000000000400ac6e01000000000000000000000000009c22000000000400de6e0100000000000000000000000000a922000000000400e66e01000000000000000000000000000000000000000400fe6e01000000000000000000000000000000000000000400fe6e01000000000000000000000000000000000000000400006f01000000000000000000000000000000000000000400046f0100000000000000000000000000b622000000000400366f0100000000000000000000000000c3220000000004003e6f01000000000000000000000000000000000000000400566f01000000000000000000000000000000000000000400566f01000000000000000000000000000000000000000400586f010000000000000000000000000000000000000004005c6f0100000000000000000000000000d0220000000004008e6f0100000000000000000000000000dd22000000000400966f01000000000000000000000000000000000000000400ae6f01000000000000000000000000000000000000000400ae6f01000000000000000000000000000000000000000400b06f01000000000000000000000000000000000000000400b46f0100000000000000000000000000ea22000000000400e66f0100000000000000000000000000f722000000000400ee6f010000000000000000000000000000000000000004000670010000000000000000000000000000000000000004000670010000000000000000000000000000000000000004000870010000000000000000000000000000000000000004000c70010000000000000000000000000004230000000004003e70010000000000000000000000000011230000000004004670010000000000000000000000000000000000000004005e70010000000000000000000000000000000000000004005e7001000000000000000000000000000000000000000400607001000000000000000000000000000000000000000400647001000000000000000000000000001e23000000000400967001000000000000000000000000002b230000000004009e7001000000000000000000000000000000000000000400b67001000000000000000000000000000000000000000400b67001000000000000000000000000000000000000000400b87001000000000000000000000000000000000000000400bc7001000000000000000000000000003823000000000400ee7001000000000000000000000000004523000000000400f670010000000000000000000000000000000000000004000e71010000000000000000000000000000000000000004000e7101000000000000000000000000000000000000000400107101000000000000000000000000000000000000000400127101000000000000000000000000005223000002000400c2cd0100000000007e00000000000000d72300000000040040710100000000000000000000000000e42300000000040048710100000000000000000000000000000000000000040060710100000000000000000000000000000000000000040060710100000000000000000000000000000000000000040062710100000000000000000000000000000000000000040066710100000000000000000000000000f12300000000040098710100000000000000000000000000fe23000000000400a07101000000000000000000000000000000000000000400b87101000000000000000000000000000000000000000400b87101000000000000000000000000000000000000000400ba7101000000000000000000000000000000000000000400bc7101000000000000000000000000000b240000020004004acd01000000000078000000000000009124000000000400ea7101000000000000000000000000009e24000000000400f271010000000000000000000000000000000000000004000a72010000000000000000000000000000000000000004000a72010000000000000000000000000000000000000004000c720100000000000000000000000000000000000000040010720100000000000000000000000000ab2400000000040036720100000000000000000000000000b8240000000004003e72010000000000000000000000000000000000000004005872010000000000000000000000000000000000000004005872010000000000000000000000000000000000000004005a72010000000000000000000000000000000000000004005e720100000000000000000000000000c52400000000040090720100000000000000000000000000d224000000000400987201000000000000000000000000000000000000000400b07201000000000000000000000000000000000000000400b07201000000000000000000000000000000000000000400b27201000000000000000000000000000000000000000400b6720100000000000000000000000000df24000000000400e8720100000000000000000000000000ec24000000000400f072010000000000000000000000000000000000000004000873010000000000000000000000000000000000000004000873010000000000000000000000000000000000000004000a730100000000000000000000000000000000000000040010730100000000000000000000000000f92400000200040086ca0100000000006200000000000000322500000200040050cb010000000000300000000000000072250000000004006e7301000000000000000000000000007f250000000004007873010000000000000000000000000000000000000004008e73010000000000000000000000000000000000000004008e7301000000000000000000000000000000000000000400907301000000000000000000000000000000000000000400947301000000000000000000000000008c25000000000400b87301000000000000000000000000009925000000000400c07301000000000000000000000000000000000000000400da7301000000000000000000000000000000000000000400da7301000000000000000000000000000000000000000400dc7301000000000000000000000000000000000000000400e0730100000000000000000000000000a62500000000040006740100000000000000000000000000b3250000000004000e74010000000000000000000000000000000000000004002874010000000000000000000000000000000000000004002874010000000000000000000000000000000000000004002a74010000000000000000000000000000000000000004002e740100000000000000000000000000c025000002000400e6cc010000000000640000000000000005260000000004008474010000000000000000000000000012260000000004008c7401000000000000000000000000001f260000000004009c7401000000000000000000000000002c26000000000400a47401000000000000000000000000000000000000000400bc7401000000000000000000000000000000000000000400bc7401000000000000000000000000000000000000000400be7401000000000000000000000000000000000000000400c27401000000000000000000000000003926000000000400187501000000000000000000000000004626000000000400207501000000000000000000000000005326000000000400307501000000000000000000000000006026000000000400387501000000000000000000000000000000000000000400507501000000000000000000000000006d260000020004005075010000000000bc0000000000000000000000000004005075010000000000000000000000000000000000000004005275010000000000000000000000000000000000000004005a750100000000000000000000000000b0260000020004000c760100000000009a00000000000000f626000002000400a676010000000000dc0000000000000000000000000004000c76010000000000000000000000000000000000000004000c76010000000000000000000000000000000000000004000e76010000000000000000000000000000000000000004001676010000000000000000000000000038270000000004002c7601000000000000000000000000004527000001000100a00201000000000040000000000000000000000000000400a67601000000000000000000000000000000000000000400a67601000000000000000000000000000000000000000400aa7601000000000000000000000000000000000000000400b676010000000000000000000000000083270000020004008277010000000000ee1a000000000000000000000000040082770100000000000000000000000000c72700000000050040c90200000000000000000000000000d12700000000050048c90200000000000000000000000000db2700000000050050c90200000000000000000000000000e52700000000050058c90200000000000000000000000000ef2700000000050060c90200000000000000000000000000f92700000000050068c90200000000000000000000000000032800000000050070c902000000000000000000000000000d2800000000050078c9020000000000000000000000000000000000000004008277010000000000000000000000000000000000000004008477010000000000000000000000000000000000000004009e77010000000000000000000000000017280000000004001e78010000000000000000000000000024280000000004003278010000000000000000000000000031280000000004007e7801000000000000000000000000003e28000000000400927801000000000000000000000000004b28000000000400dc7801000000000000000000000000005828000000000400f678010000000000000000000000000065280000000004003c7901000000000000000000000000007228000000000400527901000000000000000000000000000000000000000400709201000000000000000000000000007f280000020004007092010000000000f00000000000000000000000000004007092010000000000000000000000000000000000000004007292010000000000000000000000000000000000000004007a9201000000000000000000000000000000000000000400609301000000000000000000000000000000000000000400609301000000000000000000000000000000000000000400629301000000000000000000000000000000000000000400689301000000000000000000000000000000000000000400dc930100000000000000000000000000bd28000002000400dc9301000000000014040000000000000000000000000400dc9301000000000000000000000000000000000000000400de9301000000000000000000000000000000000000000400f8930100000000000000000000000000ff28000002000400f0970100000000003c000000000000003929000000000400be9401000000000000000000000000004729000001000100c0030100000000001c00000000000000502900000200040036980100000000004c00000000000000892900000200040082980100000000004c00000000000000d429000002000400e2bb0100000000000e00000000000000072a00000000040036970100000000000000000000000000152a0000000004004a970100000000000000000000000000232a00000000040054970100000000000000000000000000312a0000000004005e9701000000000000000000000000003e2a000000000400689701000000000000000000000000004c2a00000100010060030100000000002100000000000000552a00000000040072970100000000000000000000000000632a000001000100900301000000000024000000000000006c2a000000000400809701000000000000000000000000007a2a0000000004008a970100000000000000000000000000882a00000100010030030100000000002100000000000000912a000000000400949701000000000000000000000000009f2a0000000004009e970100000000000000000000000000ad2a000000000400a8970100000000000000000000000000bb2a00000100010000030100000000002300000000000000c42a000000000400b6970100000000000000000000000000d12a00000100010000040100000000001000000000000000fc2a000000000400d09701000000000000000000000000000a2b00000100010048040100000000001000000000000000352b0000020004002c980100000000000a000000000000006b2b000000000400e29701000000000000000000000000000000000000000400f09701000000000000000000000000000000000000000400f0970100000000000000000000000000792b00000000040008980100000000000000000000000000872b0000000004001698010000000000000000000000000000000000000004002c98010000000000000000000000000000000000000004002c980100000000000000000000000000000000000000040036980100000000000000000000000000000000000000040036980100000000000000000000000000952b00000000040054980100000000000000000000000000a32b0000000004005e980100000000000000000000000000b12b0000000004006c980100000000000000000000000000000000000000040082980100000000000000000000000000000000000000040082980100000000000000000000000000bf2b000000000400a2980100000000000000000000000000cd2b000000000400ac980100000000000000000000000000db2b000000000400c2980100000000000000000000000000e92b00000100010058040100000000000d000000000000000000000000000400ce980100000000000000000000000000142c000002000400ce98010000000000f4000000000000000000000000000400ce980100000000000000000000000000532c0000000004009a990100000000000000000000000000612c000000000400ae9901000000000000000000000000006f2c000000000400b89901000000000000000000000000000000000000000400c29901000000000000000000000000000000000000000400c29901000000000000000000000000000000000000000400c49901000000000000000000000000000000000000000400dc9901000000000000000000000000007d2c000000000400e29901000000000000000000000000008b2c000001000600e0c9020000000000a800000000000000b32c000000000400ee990100000000000000000000000000c12c000000000400989b0100000000000000000000000000cf2c000000000400da9b0100000000000000000000000000dd2c0000000004000a9d0100000000000000000000000000eb2c000000000400149d0100000000000000000000000000f92c000000000400229d0100000000000000000000000000072d000000000400369d0100000000000000000000000000152d000000000400409d0100000000000000000000000000232d000000000400549d0100000000000000000000000000312d0000000004005c9d01000000000000000000000000003f2d000001000100e0020100000000002000000000000000692d000000000400669d0100000000000000000000000000772d0000000004006e9d0100000000000000000000000000852d000000000400789d0100000000000000000000000000932d000000000400809d01000000000000000000000000000000000000000400969d01000000000000000000000000000000000000000400969d01000000000000000000000000000000000000000400989d01000000000000000000000000000000000000000400b29d0100000000000000000000000000a12d000000000400b29d0100000000000000000000000000af2d000000000400d09d0100000000000000000000000000bd2d0000000004001c9e0100000000000000000000000000cb2d000000000400c49e0100000000000000000000000000d92d00000000040014a10100000000000000000000000000e72d0000000004001ea10100000000000000000000000000f52d0000000004002ca10100000000000000000000000000032e00000000040040a10100000000000000000000000000112e00000000040058a101000000000000000000000000001f2e00000000040060a101000000000000000000000000002d2e0000000004006aa101000000000000000000000000003b2e00000000040072a10100000000000000000000000000000000000000040088a10100000000000000000000000000000000000000040088a1010000000000000000000000000000000000000004008aa10100000000000000000000000000000000000000040098a10100000000000000000000000000492e0000020004005ea20100000000005200000000000000912e000002000400b0a20100000000003400000000000000eb2e0000000004003ca20100000000000000000000000000f92e0000010001007004010000000000190000000000000000000000000004005ea2010000000000000000000000000000000000000004005ea20100000000000000000000000000000000000000040060a20100000000000000000000000000000000000000040066a201000000000000000000000000000000000000000400b0a201000000000000000000000000000000000000000400b0a201000000000000000000000000000000000000000400b2a201000000000000000000000000000000000000000400b4a20100000000000000000000000000022f000002000400e4a201000000000074000000000000000000000000000400e4a201000000000000000000000000000000000000000400e4a201000000000000000000000000000000000000000400e6a201000000000000000000000000000000000000000400eca201000000000000000000000000004d2f000002000400b2c50100000000006200000000000000000000000000040058a30100000000000000000000000000802f00000200040058a30100000000003600000000000000000000000000040058a3010000000000000000000000000000000000000004005aa3010000000000000000000000000000000000000004005ca3010000000000000000000000000000000000000004008ea3010000000000000000000000000000000000000004008ea30100000000000000000000000000000000000000040090a3010000000000000000000000000000000000000004009ca301000000000000000000000000000000000000000400faa301000000000000000000000000000000000000000400faa3010000000000000000000000000000000000000004001ca4010000000000000000000000000000000000000004001ca4010000000000000000000000000000000000000004001ea40100000000000000000000000000000000000000040024a40100000000000000000000000000000000000000040056a40100000000000000000000000000000000000000040056a40100000000000000000000000000000000000000040058a40100000000000000000000000000000000000000040066a40100000000000000000000000000cd2f00000000040082a40100000000000000000000000000db2f000001000100c2040100000000000b000000000000000730000000000400dea40100000000000000000000000000153000000000040038a50100000000000000000000000000000000000000040052a50100000000000000000000000000000000000000040052a50100000000000000000000000000000000000000040094a50100000000000000000000000000233000000200040094a50100000000005000000000000000000000000000040094a50100000000000000000000000000000000000000040096a501000000000000000000000000000000000000000400a2a501000000000000000000000000000000000000000400e4a501000000000000000000000000000631000002000400e4a501000000000074000000000000000000000000000400e4a501000000000000000000000000000000000000000400e6a501000000000000000000000000000000000000000400eea50100000000000000000000000000da31000002000400e2c40100000000005200000000000000863200000000040044a60100000000000000000000000000943200000100010090040100000000001c00000000000000000000000000040058a60100000000000000000000000000000000000000040058a6010000000000000000000000000000000000000004005aa60100000000000000000000000000000000000000040066a601000000000000000000000000000000000000000400bca601000000000000000000000000009d32000002000400bca601000000000082000000000000000000000000000400bca601000000000000000000000000000000000000000400bea601000000000000000000000000000000000000000400c6a6010000000000000000000000000000000000000004003ea7010000000000000000000000000025330000020004003ea7010000000000960100000000000000000000000004003ea70100000000000000000000000000000000000000040040a70100000000000000000000000000000000000000040054a70100000000000000000000000000af33000000000400aca80100000000000000000000000000bd33000000000400b6a80100000000000000000000000000cb33000000000400c0a801000000000000000000000000000000000000000400d4a801000000000000000000000000000000000000000400d4a80100000000000000000000000000000000000000040046a90100000000000000000000000000d93300000200040046a90100000000009200000000000000000000000000040046a90100000000000000000000000000000000000000040048a9010000000000000000000000000000000000000004004aa9010000000000000000000000000034340000000004004ea901000000000000000000000000004234000000000100600101000000000000000000000000004c340000000004005ca90100000000000000000000000000553400000000040062a9010000000000000000000000000063340000010001009b050100000000000f000000000000008e340000000004006ea90100000000000000000000000000973400000000040074a90100000000000000000000000000a53400000100010090050100000000000b00000000000000d03400000000040080a90100000000000000000000000000d93400000000040084a90100000000000000000000000000e73400000100010060050100000000000f0000000000000012350000000004008ca901000000000000000000000000002035000001000100700501000000000020000000000000004b3500000000040098a9010000000000000000000000000054350000000004009ea901000000000000000000000000006235000000000400aea901000000000000000000000000006b35000000000400b2a9010000000000000000000000000079350000010001001d050100000000000700000000000000a435000000000400baa90100000000000000000000000000b23500000100010028050100000000002000000000000000dd3500000200040030c201000000000098000000000000000000000000000400d8a901000000000000000000000000002336000002000400d8a901000000000002000000000000000000000000000400d8a901000000000000000000000000000000000000000400daa901000000000000000000000000000000000000000400daa90100000000000000000000000000000000000000040010aa0100000000000000000000000000000000000000040010aa0100000000000000000000000000000000000000040014aa0100000000000000000000000000000000000000040038aa0100000000000000000000000000623600000000040032ab01000000000000000000000000007036000001000100fd040100000000000f000000000000000000000000000400d0ab01000000000000000000000000009c36000002000400d0ab0100000000007a000000000000000000000000000400d0ab01000000000000000000000000000000000000000400d2ab01000000000000000000000000000000000000000400d6ab010000000000000000000000000000000000000004004aac010000000000000000000000000000000000000004004aac010000000000000000000000000000000000000004004cac0100000000000000000000000000000000000000040050ac01000000000000000000000000000000000000000400ccac0100000000000000000000000000dd36000002000400ccac01000000000060010000000000000000000000000400ccac01000000000000000000000000000000000000000400d0ac01000000000000000000000000000000000000000400f4ac010000000000000000000000000000000000000004002cae010000000000000000000000000000000000000004002cae0100000000000000000000000000000000000000040030ae0100000000000000000000000000000000000000040060ae0100000000000000000000000000193700000000040052af01000000000000000000000000002737000001000100f1040100000000000c00000000000000533700000000040096af01000000000000000000000000006137000000000400b2af01000000000000000000000000006f370000000004005cb001000000000000000000000000007d370000000004008ab001000000000000000000000000008b37000000000400f0b00100000000000000000000000000993700000000040080b10100000000000000000000000000a737000000000400aab10100000000000000000000000000b53700000000040072b20100000000000000000000000000c337000001000100b6040100000000000c00000000000000ee3700000000040092b20100000000000000000000000000fc37000001000100ac040100000000000a000000000000000000000000000400eeb201000000000000000000000000000000000000000400eeb20100000000000000000000000000000000000000040006b30100000000000000000000000000000000000000040006b30100000000000000000000000000000000000000040008b3010000000000000000000000000000000000000004002ab3010000000000000000000000000027380000020004002ab3010000000000040000000000000000000000000004002ab3010000000000000000000000000000000000000004002ab3010000000000000000000000000000000000000004002ab3010000000000000000000000000000000000000004002ab3010000000000000000000000000000000000000004002cb3010000000000000000000000000000000000000004002cb3010000000000000000000000000000000000000004002eb3010000000000000000000000000000000000000004002eb3010000000000000000000000000000000000000004002eb3010000000000000000000000000062380000020004002eb3010000000000020000000000000000000000000004002eb3010000000000000000000000000000000000000004002eb3010000000000000000000000000000000000000004002eb3010000000000000000000000000000000000000004002eb30100000000000000000000000000000000000000040030b30100000000000000000000000000000000000000040030b30100000000000000000000000000ec3800000000050080c90200000000000000000000000000f63800000200040030b30100000000004201000000000000000000000000040030b30100000000000000000000000000000000000000040030b30100000000000000000000000000000000000000040030b30100000000000000000000000000000000000000040032b30100000000000000000000000000000000000000040034b30100000000000000000000000000000000000000040036b30100000000000000000000000000273900000000040042b3010000000000000000000000000035390000010001003006010000000000c80000000000000000000000000004004eb30100000000000000000000000000000000000000040052b30100000000000000000000000000613900000000040056b30100000000000000000000000000000000000000040076b30100000000000000000000000000000000000000040078b30100000000000000000000000000000000000000040086b301000000000000000000000000000000000000000400a0b301000000000000000000000000000000000000000400a0b301000000000000000000000000000000000000000400a2b301000000000000000000000000000000000000000400a2b301000000000000000000000000000000000000000400a6b301000000000000000000000000000000000000000400a6b301000000000000000000000000000000000000000400aab301000000000000000000000000000000000000000400aab301000000000000000000000000000000000000000400b2b301000000000000000000000000000000000000000400b2b301000000000000000000000000000000000000000400b4b301000000000000000000000000000000000000000400b4b301000000000000000000000000000000000000000400bcb301000000000000000000000000000000000000000400bcb301000000000000000000000000000000000000000400beb301000000000000000000000000000000000000000400beb301000000000000000000000000000000000000000400c2b301000000000000000000000000000000000000000400c2b301000000000000000000000000000000000000000400cab301000000000000000000000000000000000000000400cab301000000000000000000000000000000000000000400d0b301000000000000000000000000000000000000000400d4b301000000000000000000000000000000000000000400d8b301000000000000000000000000000000000000000400f4b301000000000000000000000000000000000000000400f8b301000000000000000000000000000000000000000400fab301000000000000000000000000000000000000000400fab301000000000000000000000000000000000000000400fcb301000000000000000000000000000000000000000400fcb30100000000000000000000000000000000000000040008b40100000000000000000000000000000000000000040008b4010000000000000000000000000000000000000004000ab4010000000000000000000000000000000000000004000ab40100000000000000000000000000000000000000040014b40100000000000000000000000000000000000000040014b40100000000000000000000000000000000000000040016b4010000000000000000000000000000000000000004001ab40100000000000000000000000000000000000000040022b40100000000000000000000000000000000000000040022b40100000000000000000000000000000000000000040024b40100000000000000000000000000000000000000040024b4010000000000000000000000000000000000000004002eb40100000000000000000000000000000000000000040030b40100000000000000000000000000000000000000040034b40100000000000000000000000000000000000000040034b40100000000000000000000000000000000000000040036b40100000000000000000000000000000000000000040036b40100000000000000000000000000000000000000040042b40100000000000000000000000000000000000000040042b40100000000000000000000000000000000000000040044b40100000000000000000000000000000000000000040044b4010000000000000000000000000000000000000004004cb4010000000000000000000000000000000000000004004cb40100000000000000000000000000000000000000040050b40100000000000000000000000000000000000000040050b40100000000000000000000000000000000000000040056b40100000000000000000000000000000000000000040056b401000000000000000000000000006f3900000000040058b401000000000000000000000000007d39000001000100300a0100000000000000000000000000000000000000040058b40100000000000000000000000000a83900000200040072b4010000000000e40100000000000000000000000004006cb4010000000000000000000000000000000000000004006eb40100000000000000000000000000000000000000040072b40100000000000000000000000000000000000000040072b40100000000000000000000000000000000000000040072b40100000000000000000000000000000000000000040072b40100000000000000000000000000000000000000040072b40100000000000000000000000000000000000000040074b4010000000000000000000000000000000000000004008eb40100000000000000000000000000000000000000040090b40100000000000000000000000000000000000000040090b4010000000000000000000000000000000000000004009cb4010000000000000000000000000000000000000004009cb401000000000000000000000000000000000000000400a8b401000000000000000000000000000000000000000400acb401000000000000000000000000000000000000000400acb401000000000000000000000000000000000000000400b0b401000000000000000000000000000000000000000400b0b401000000000000000000000000000000000000000400b2b401000000000000000000000000000000000000000400b4b401000000000000000000000000000000000000000400b6b401000000000000000000000000000000000000000400b8b401000000000000000000000000000000000000000400bcb401000000000000000000000000000000000000000400beb401000000000000000000000000000000000000000400beb401000000000000000000000000000000000000000400c2b401000000000000000000000000000000000000000400c2b401000000000000000000000000000000000000000400c6b401000000000000000000000000000000000000000400cab401000000000000000000000000000000000000000400cab401000000000000000000000000000000000000000400ccb401000000000000000000000000000000000000000400ccb401000000000000000000000000000000000000000400d4b401000000000000000000000000000000000000000400d4b401000000000000000000000000000000000000000400d6b401000000000000000000000000000000000000000400d6b401000000000000000000000000000000000000000400d8b401000000000000000000000000000000000000000400d8b401000000000000000000000000000000000000000400dab401000000000000000000000000000000000000000400dab401000000000000000000000000000000000000000400dcb401000000000000000000000000000000000000000400deb401000000000000000000000000000000000000000400e0b401000000000000000000000000000000000000000400e4b401000000000000000000000000000000000000000400e8b401000000000000000000000000000000000000000400e8b401000000000000000000000000000000000000000400eab401000000000000000000000000000000000000000400eab401000000000000000000000000000000000000000400ecb401000000000000000000000000000000000000000400ecb401000000000000000000000000000000000000000400f2b401000000000000000000000000000000000000000400f2b401000000000000000000000000000000000000000400f6b401000000000000000000000000000000000000000400f6b401000000000000000000000000000000000000000400fcb401000000000000000000000000000000000000000400fcb40100000000000000000000000000e13900000200040056b6010000000000560000000000000000000000000004001cb50100000000000000000000000000000000000000040038b5010000000000000000000000000000000000000004003cb50100000000000000000000000000000000000000040062b50100000000000000000000000000000000000000040062b50100000000000000000000000000000000000000040068b50100000000000000000000000000000000000000040068b5010000000000000000000000000000000000000004006cb5010000000000000000000000000000000000000004006cb50100000000000000000000000000000000000000040076b50100000000000000000000000000000000000000040076b5010000000000000000000000000000000000000004007ab5010000000000000000000000000000000000000004007ab5010000000000000000000000000000000000000004007eb5010000000000000000000000000000000000000004007eb50100000000000000000000000000000000000000040092b50100000000000000000000000000000000000000040094b50100000000000000000000000000000000000000040094b5010000000000000000000000000000000000000004009ab5010000000000000000000000000000000000000004009ab5010000000000000000000000000000000000000004009eb5010000000000000000000000000000000000000004009eb501000000000000000000000000000000000000000400aeb501000000000000000000000000000000000000000400aeb501000000000000000000000000000000000000000400b0b501000000000000000000000000000000000000000400b0b501000000000000000000000000000000000000000400b4b501000000000000000000000000000000000000000400b8b501000000000000000000000000000000000000000400bab501000000000000000000000000000000000000000400c0b501000000000000000000000000000000000000000400ccb501000000000000000000000000000000000000000400d0b501000000000000000000000000000000000000000400d0b501000000000000000000000000000000000000000400d2b501000000000000000000000000000000000000000400d2b501000000000000000000000000000000000000000400d4b501000000000000000000000000000000000000000400d4b501000000000000000000000000000000000000000400e0b501000000000000000000000000000000000000000400e0b501000000000000000000000000000000000000000400eab501000000000000000000000000000000000000000400eeb50100000000000000000000000000000000000000040002b60100000000000000000000000000000000000000040010b60100000000000000000000000000000000000000040010b60100000000000000000000000000000000000000040018b60100000000000000000000000000000000000000040018b60100000000000000000000000000000000000000040020b60100000000000000000000000000000000000000040020b60100000000000000000000000000000000000000040030b60100000000000000000000000000000000000000040030b60100000000000000000000000000000000000000040040b60100000000000000000000000000000000000000040042b60100000000000000000000000000000000000000040046b6010000000000000000000000000000000000000004004eb60100000000000000000000000000000000000000040050b60100000000000000000000000000000000000000040050b60100000000000000000000000000000000000000040056b60100000000000000000000000000000000000000040056b60100000000000000000000000000000000000000040056b60100000000000000000000000000000000000000040056b60100000000000000000000000000000000000000040056b60100000000000000000000000000000000000000040056b60100000000000000000000000000000000000000040058b60100000000000000000000000000000000000000040062b60100000000000000000000000000000000000000040072b60100000000000000000000000000000000000000040076b60100000000000000000000000000000000000000040084b60100000000000000000000000000000000000000040086b60100000000000000000000000000000000000000040098b6010000000000000000000000000000000000000004009cb6010000000000000000000000000000000000000004009eb601000000000000000000000000000000000000000400a8b601000000000000000000000000000000000000000400acb601000000000000000000000000000000000000000400acb60100000000000000000000000000283a00000000050088c90200000000000000000000000000323a00000000050090c902000000000000000000000000003c3a000002000400acb601000000000078030000000000000000000000000400acb601000000000000000000000000000000000000000400acb601000000000000000000000000000000000000000400acb601000000000000000000000000000000000000000400aeb601000000000000000000000000000000000000000400aeb601000000000000000000000000000000000000000400aeb601000000000000000000000000000000000000000400c0b601000000000000000000000000000000000000000400c4b601000000000000000000000000000000000000000400c4b601000000000000000000000000000000000000000400c6b601000000000000000000000000000000000000000400c6b601000000000000000000000000000000000000000400ceb601000000000000000000000000000000000000000400ceb601000000000000000000000000000000000000000400d2b601000000000000000000000000000000000000000400d6b601000000000000000000000000000000000000000400dab601000000000000000000000000000000000000000400dab601000000000000000000000000000000000000000400deb601000000000000000000000000000000000000000400deb601000000000000000000000000000000000000000400f0b601000000000000000000000000000000000000000400f0b601000000000000000000000000000000000000000400f4b601000000000000000000000000000000000000000400f4b601000000000000000000000000000000000000000400f6b601000000000000000000000000000000000000000400fab601000000000000000000000000000000000000000400fab601000000000000000000000000000000000000000400feb601000000000000000000000000000000000000000400feb60100000000000000000000000000000000000000040000b70100000000000000000000000000000000000000040000b70100000000000000000000000000000000000000040002b70100000000000000000000000000000000000000040002b70100000000000000000000000000000000000000040006b70100000000000000000000000000000000000000040006b7010000000000000000000000000000000000000004000eb70100000000000000000000000000000000000000040012b70100000000000000000000000000000000000000040016b70100000000000000000000000000000000000000040016b7010000000000000000000000000000000000000004001ab7010000000000000000000000000000000000000004001ab7010000000000000000000000000000000000000004001eb7010000000000000000000000000000000000000004001eb70100000000000000000000000000000000000000040022b70100000000000000000000000000000000000000040026b70100000000000000000000000000000000000000040026b70100000000000000000000000000000000000000040028b7010000000000000000000000000000000000000004002cb70100000000000000000000000000000000000000040030b70100000000000000000000000000000000000000040030b70100000000000000000000000000000000000000040034b70100000000000000000000000000000000000000040038b7010000000000000000000000000000000000000004003cb7010000000000000000000000000000000000000004003cb7010000000000000000000000000000000000000004003eb70100000000000000000000000000000000000000040042b70100000000000000000000000000000000000000040046b70100000000000000000000000000000000000000040046b70100000000000000000000000000000000000000040048b70100000000000000000000000000000000000000040048b7010000000000000000000000000000000000000004004cb7010000000000000000000000000000000000000004004cb7010000000000000000000000000000000000000004006ab7010000000000000000000000000000000000000004006ab7010000000000000000000000000000000000000004006eb7010000000000000000000000000000000000000004006eb70100000000000000000000000000000000000000040072b70100000000000000000000000000000000000000040076b7010000000000000000000000000000000000000004007eb70100000000000000000000000000000000000000040082b70100000000000000000000000000000000000000040086b7010000000000000000000000000000000000000004008ab7010000000000000000000000000000000000000004008eb70100000000000000000000000000000000000000040092b70100000000000000000000000000000000000000040092b70100000000000000000000000000000000000000040096b70100000000000000000000000000000000000000040096b7010000000000000000000000000000000000000004009ab7010000000000000000000000000000000000000004009ab7010000000000000000000000000000000000000004009eb701000000000000000000000000000000000000000400a2b701000000000000000000000000000000000000000400a2b701000000000000000000000000000000000000000400a8b701000000000000000000000000000000000000000400acb701000000000000000000000000000000000000000400aeb701000000000000000000000000000000000000000400aeb701000000000000000000000000000000000000000400b4b701000000000000000000000000000000000000000400b4b701000000000000000000000000000000000000000400b8b701000000000000000000000000000000000000000400b8b701000000000000000000000000000000000000000400bab701000000000000000000000000000000000000000400beb701000000000000000000000000000000000000000400beb701000000000000000000000000000000000000000400c2b701000000000000000000000000000000000000000400c2b701000000000000000000000000000000000000000400cab701000000000000000000000000000000000000000400cab701000000000000000000000000000000000000000400ceb701000000000000000000000000000000000000000400ceb701000000000000000000000000000000000000000400d0b701000000000000000000000000000000000000000400d0b701000000000000000000000000000000000000000400d4b701000000000000000000000000000000000000000400d4b701000000000000000000000000000000000000000400d8b701000000000000000000000000000000000000000400d8b701000000000000000000000000000000000000000400dab701000000000000000000000000000000000000000400dab701000000000000000000000000000000000000000400dcb701000000000000000000000000000000000000000400dcb701000000000000000000000000000000000000000400e0b701000000000000000000000000000000000000000400e4b701000000000000000000000000000000000000000400ecb701000000000000000000000000000000000000000400ecb701000000000000000000000000000000000000000400f0b701000000000000000000000000000000000000000400f2b701000000000000000000000000000000000000000400f2b701000000000000000000000000000000000000000400f6b701000000000000000000000000000000000000000400f6b701000000000000000000000000000000000000000400fab701000000000000000000000000000000000000000400feb701000000000000000000000000000000000000000400feb70100000000000000000000000000000000000000040000b80100000000000000000000000000000000000000040000b80100000000000000000000000000000000000000040008b80100000000000000000000000000000000000000040008b8010000000000000000000000000000000000000004000ab8010000000000000000000000000000000000000004000ab8010000000000000000000000000000000000000004000cb8010000000000000000000000000000000000000004000cb80100000000000000000000000000000000000000040010b80100000000000000000000000000000000000000040010b80100000000000000000000000000000000000000040016b80100000000000000000000000000000000000000040016b8010000000000000000000000000000000000000004001eb8010000000000000000000000000000000000000004001eb80100000000000000000000000000000000000000040024b80100000000000000000000000000000000000000040024b80100000000000000000000000000000000000000040028b80100000000000000000000000000000000000000040028b8010000000000000000000000000000000000000004002ab8010000000000000000000000000000000000000004002eb8010000000000000000000000000000000000000004002eb80100000000000000000000000000000000000000040030b80100000000000000000000000000000000000000040030b80100000000000000000000000000000000000000040038b80100000000000000000000000000000000000000040038b8010000000000000000000000000000000000000004003ab8010000000000000000000000000000000000000004003ab8010000000000000000000000000000000000000004003cb8010000000000000000000000000000000000000004003cb8010000000000000000000000000000000000000004003eb8010000000000000000000000000000000000000004003eb80100000000000000000000000000000000000000040040b80100000000000000000000000000000000000000040040b80100000000000000000000000000000000000000040042b80100000000000000000000000000000000000000040042b80100000000000000000000000000000000000000040048b8010000000000000000000000000000000000000004004cb8010000000000000000000000000000000000000004004cb8010000000000000000000000000000000000000004004eb8010000000000000000000000000000000000000004004eb80100000000000000000000000000000000000000040056b80100000000000000000000000000000000000000040056b80100000000000000000000000000000000000000040058b80100000000000000000000000000000000000000040058b8010000000000000000000000000000000000000004005ab8010000000000000000000000000000000000000004005ab8010000000000000000000000000000000000000004005cb8010000000000000000000000000000000000000004005cb801000000000000000000000000006b3a00000000040060b80100000000000000000000000000793a00000000040068b8010000000000000000000000000000000000000004007eb80100000000000000000000000000000000000000040084b80100000000000000000000000000000000000000040092b80100000000000000000000000000000000000000040092b80100000000000000000000000000000000000000040096b80100000000000000000000000000000000000000040098b8010000000000000000000000000000000000000004009cb8010000000000000000000000000000000000000004009eb8010000000000000000000000000000000000000004009eb801000000000000000000000000000000000000000400a2b801000000000000000000000000000000000000000400a2b801000000000000000000000000000000000000000400a4b801000000000000000000000000000000000000000400a4b801000000000000000000000000000000000000000400a6b801000000000000000000000000000000000000000400a8b801000000000000000000000000000000000000000400a8b801000000000000000000000000000000000000000400aab801000000000000000000000000000000000000000400b4b801000000000000000000000000000000000000000400b8b801000000000000000000000000000000000000000400bcb801000000000000000000000000000000000000000400bcb801000000000000000000000000000000000000000400c0b801000000000000000000000000000000000000000400c0b801000000000000000000000000000000000000000400c6b801000000000000000000000000000000000000000400c6b801000000000000000000000000000000000000000400c8b801000000000000000000000000000000000000000400c8b801000000000000000000000000000000000000000400ccb801000000000000000000000000000000000000000400ceb801000000000000000000000000000000000000000400d0b801000000000000000000000000000000000000000400d0b801000000000000000000000000000000000000000400d4b801000000000000000000000000000000000000000400d6b801000000000000000000000000000000000000000400d8b801000000000000000000000000000000000000000400d8b801000000000000000000000000000000000000000400dab801000000000000000000000000000000000000000400dab801000000000000000000000000000000000000000400deb801000000000000000000000000000000000000000400deb801000000000000000000000000000000000000000400e0b801000000000000000000000000000000000000000400e0b801000000000000000000000000000000000000000400e4b801000000000000000000000000000000000000000400e6b801000000000000000000000000000000000000000400e6b801000000000000000000000000000000000000000400e8b801000000000000000000000000000000000000000400e8b801000000000000000000000000000000000000000400eab801000000000000000000000000000000000000000400eeb801000000000000000000000000000000000000000400f2b801000000000000000000000000000000000000000400f4b801000000000000000000000000000000000000000400f6b801000000000000000000000000000000000000000400f8b801000000000000000000000000000000000000000400f8b801000000000000000000000000000000000000000400fab801000000000000000000000000000000000000000400fab801000000000000000000000000000000000000000400fcb801000000000000000000000000000000000000000400fcb80100000000000000000000000000000000000000040000b90100000000000000000000000000000000000000040000b90100000000000000000000000000000000000000040004b90100000000000000000000000000000000000000040006b90100000000000000000000000000000000000000040008b9010000000000000000000000000000000000000004000cb9010000000000000000000000000000000000000004000cb90100000000000000000000000000000000000000040010b90100000000000000000000000000000000000000040010b90100000000000000000000000000000000000000040012b90100000000000000000000000000000000000000040012b90100000000000000000000000000000000000000040018b90100000000000000000000000000000000000000040018b9010000000000000000000000000000000000000004001cb90100000000000000000000000000000000000000040020b90100000000000000000000000000000000000000040024b9010000000000000000000000000000000000000004002ab90100000000000000000000000000000000000000040030b90100000000000000000000000000000000000000040030b90100000000000000000000000000000000000000040032b90100000000000000000000000000000000000000040032b90100000000000000000000000000000000000000040034b90100000000000000000000000000000000000000040034b90100000000000000000000000000000000000000040038b9010000000000000000000000000000000000000004003ab9010000000000000000000000000000000000000004003cb90100000000000000000000000000000000000000040040b90100000000000000000000000000000000000000040040b90100000000000000000000000000000000000000040042b90100000000000000000000000000000000000000040042b90100000000000000000000000000000000000000040044b90100000000000000000000000000000000000000040044b90100000000000000000000000000000000000000040048b90100000000000000000000000000000000000000040048b9010000000000000000000000000000000000000004004ab9010000000000000000000000000000000000000004004ab9010000000000000000000000000000000000000004004eb90100000000000000000000000000000000000000040050b90100000000000000000000000000000000000000040054b90100000000000000000000000000000000000000040056b90100000000000000000000000000000000000000040056b9010000000000000000000000000000000000000004005ab9010000000000000000000000000000000000000004005ab9010000000000000000000000000000000000000004005cb9010000000000000000000000000000000000000004005cb9010000000000000000000000000000000000000004005eb9010000000000000000000000000000000000000004005eb90100000000000000000000000000000000000000040062b90100000000000000000000000000000000000000040062b90100000000000000000000000000000000000000040068b90100000000000000000000000000000000000000040068b9010000000000000000000000000000000000000004006cb9010000000000000000000000000000000000000004006cb90100000000000000000000000000000000000000040072b90100000000000000000000000000000000000000040072b90100000000000000000000000000000000000000040098b90100000000000000000000000000000000000000040098b9010000000000000000000000000000000000000004009cb901000000000000000000000000000000000000000400a0b901000000000000000000000000000000000000000400a2b901000000000000000000000000000000000000000400a8b901000000000000000000000000000000000000000400b6b901000000000000000000000000000000000000000400bab901000000000000000000000000000000000000000400bab901000000000000000000000000000000000000000400bcb901000000000000000000000000000000000000000400bcb901000000000000000000000000000000000000000400beb901000000000000000000000000000000000000000400beb901000000000000000000000000000000000000000400cab901000000000000000000000000000000000000000400cab901000000000000000000000000000000000000000400d4b901000000000000000000000000000000000000000400d8b901000000000000000000000000000000000000000400e6b901000000000000000000000000000000000000000400e6b901000000000000000000000000000000000000000400eeb901000000000000000000000000000000000000000400eeb901000000000000000000000000000000000000000400f2b901000000000000000000000000000000000000000400f2b901000000000000000000000000000000000000000400f6b901000000000000000000000000000000000000000400f6b90100000000000000000000000000000000000000040006ba0100000000000000000000000000000000000000040008ba0100000000000000000000000000000000000000040008ba010000000000000000000000000000000000000004000cba010000000000000000000000000000000000000004000cba0100000000000000000000000000000000000000040020ba0100000000000000000000000000000000000000040024ba0100000000000000000000000000000000000000040024ba0100000000000000000000000000000000000000040024ba0100000000000000000000000000000000000000040024ba0100000000000000000000000000000000000000040024ba0100000000000000000000000000000000000000040026ba0100000000000000000000000000000000000000040026ba0100000000000000000000000000000000000000040028ba0100000000000000000000000000000000000000040032ba0100000000000000000000000000000000000000040032ba0100000000000000000000000000873a00000200040032ba0100000000007e01000000000000000000000000040032ba0100000000000000000000000000000000000000040032ba0100000000000000000000000000000000000000040032ba0100000000000000000000000000000000000000040034ba0100000000000000000000000000000000000000040044ba010000000000000000000000000000000000000004004aba010000000000000000000000000000000000000004004aba0100000000000000000000000000000000000000040052ba0100000000000000000000000000000000000000040052ba0100000000000000000000000000000000000000040056ba0100000000000000000000000000000000000000040056ba010000000000000000000000000000000000000004005eba010000000000000000000000000000000000000004005eba0100000000000000000000000000000000000000040060ba0100000000000000000000000000000000000000040064ba0100000000000000000000000000000000000000040064ba0100000000000000000000000000000000000000040068ba010000000000000000000000000000000000000004006cba0100000000000000000000000000ae3a00000000040086ba010000000000000000000000000000000000000004008eba010000000000000000000000000000000000000004008eba0100000000000000000000000000000000000000040090ba0100000000000000000000000000000000000000040092ba0100000000000000000000000000000000000000040096ba010000000000000000000000000000000000000004009aba01000000000000000000000000000000000000000400a0ba01000000000000000000000000000000000000000400a0ba01000000000000000000000000000000000000000400a2ba01000000000000000000000000000000000000000400a4ba01000000000000000000000000000000000000000400a8ba01000000000000000000000000000000000000000400acba01000000000000000000000000000000000000000400aeba01000000000000000000000000000000000000000400aeba01000000000000000000000000000000000000000400b2ba01000000000000000000000000000000000000000400b2ba01000000000000000000000000000000000000000400b4ba01000000000000000000000000000000000000000400baba01000000000000000000000000000000000000000400baba01000000000000000000000000000000000000000400c0ba01000000000000000000000000000000000000000400c0ba01000000000000000000000000000000000000000400caba01000000000000000000000000000000000000000400ceba01000000000000000000000000000000000000000400d0ba01000000000000000000000000000000000000000400d2ba01000000000000000000000000000000000000000400d2ba01000000000000000000000000000000000000000400d4ba01000000000000000000000000000000000000000400d8ba01000000000000000000000000000000000000000400e0ba01000000000000000000000000000000000000000400e0ba01000000000000000000000000000000000000000400e6ba01000000000000000000000000000000000000000400e6ba01000000000000000000000000000000000000000400f0ba01000000000000000000000000000000000000000400f4ba01000000000000000000000000000000000000000400f6ba01000000000000000000000000000000000000000400f8ba01000000000000000000000000000000000000000400f8ba01000000000000000000000000000000000000000400faba01000000000000000000000000000000000000000400feba0100000000000000000000000000000000000000040000bb0100000000000000000000000000000000000000040000bb0100000000000000000000000000000000000000040004bb0100000000000000000000000000000000000000040004bb0100000000000000000000000000000000000000040006bb0100000000000000000000000000000000000000040008bb010000000000000000000000000000000000000004000cbb010000000000000000000000000000000000000004000cbb010000000000000000000000000000000000000004000ebb010000000000000000000000000000000000000004000ebb010000000000000000000000000000000000000004001ebb010000000000000000000000000000000000000004001ebb0100000000000000000000000000000000000000040022bb0100000000000000000000000000000000000000040022bb0100000000000000000000000000000000000000040026bb010000000000000000000000000000000000000004002ebb0100000000000000000000000000000000000000040040bb0100000000000000000000000000000000000000040040bb0100000000000000000000000000000000000000040042bb0100000000000000000000000000000000000000040044bb0100000000000000000000000000000000000000040048bb010000000000000000000000000000000000000004004cbb0100000000000000000000000000000000000000040052bb0100000000000000000000000000000000000000040052bb0100000000000000000000000000000000000000040054bb0100000000000000000000000000000000000000040058bb010000000000000000000000000000000000000004005cbb010000000000000000000000000000000000000004005cbb010000000000000000000000000000000000000004005ebb010000000000000000000000000000000000000004005ebb0100000000000000000000000000000000000000040068bb0100000000000000000000000000000000000000040068bb010000000000000000000000000000000000000004006cbb010000000000000000000000000000000000000004006cbb0100000000000000000000000000000000000000040072bb0100000000000000000000000000000000000000040072bb0100000000000000000000000000000000000000040074bb0100000000000000000000000000000000000000040078bb0100000000000000000000000000000000000000040078bb010000000000000000000000000000000000000004007cbb010000000000000000000000000000000000000004007cbb0100000000000000000000000000000000000000040080bb0100000000000000000000000000000000000000040080bb0100000000000000000000000000000000000000040084bb0100000000000000000000000000000000000000040084bb0100000000000000000000000000000000000000040088bb0100000000000000000000000000000000000000040090bb0100000000000000000000000000000000000000040096bb010000000000000000000000000000000000000004009cbb01000000000000000000000000000000000000000400acbb01000000000000000000000000000000000000000400b0bb01000000000000000000000000000000000000000400b0bb0100000000000000000000000000bc3a000002000400b0bb01000000000012000000000000000000000000000400b0bb01000000000000000000000000000000000000000400b0bb01000000000000000000000000000000000000000400b0bb01000000000000000000000000000000000000000400b0bb0100000000000000000000000000163b000000000400b6bb0100000000000000000000000000243b000001000100cd050100000000000b000000000000000000000000000400c2bb01000000000000000000000000000000000000000400c2bb01000000000000000000000000000000000000000400c2bb0100000000000000000000000000503b000002000400c2bb01000000000012000000000000000000000000000400c2bb01000000000000000000000000000000000000000400c2bb01000000000000000000000000000000000000000400c2bb01000000000000000000000000000000000000000400c2bb0100000000000000000000000000ad3b000000000400c8bb0100000000000000000000000000bb3b000001000100d8050100000000000e000000000000000000000000000400d4bb01000000000000000000000000000000000000000400d4bb01000000000000000000000000000000000000000400d4bb01000000000000000000000000000000000000000400d4bb01000000000000000000000000000000000000000400d4bb01000000000000000000000000000000000000000400d4bb01000000000000000000000000000000000000000400d6bb01000000000000000000000000000000000000000400d6bb01000000000000000000000000000000000000000400d8bb01000000000000000000000000000000000000000400e2bb01000000000000000000000000000000000000000400e2bb01000000000000000000000000000000000000000400e2bb01000000000000000000000000000000000000000400e2bb01000000000000000000000000000000000000000400e2bb01000000000000000000000000000000000000000400e4bb01000000000000000000000000000000000000000400e4bb01000000000000000000000000000000000000000400e4bb01000000000000000000000000000000000000000400e6bb01000000000000000000000000000000000000000400f0bb01000000000000000000000000000000000000000400f0bb01000000000000000000000000000000000000000400f0bb01000000000000000000000000000000000000000400f0bb01000000000000000000000000000000000000000400f0bb01000000000000000000000000000000000000000400f0bb01000000000000000000000000000000000000000400f2bb01000000000000000000000000000000000000000400f2bb01000000000000000000000000000000000000000400f4bb01000000000000000000000000000000000000000400febb01000000000000000000000000000000000000000400febb0100000000000000000000000000e73b000002000400febb01000000000070000000000000000000000000000400febb01000000000000000000000000000000000000000400febb01000000000000000000000000000000000000000400febb0100000000000000000000000000000000000000040000bc0100000000000000000000000000000000000000040002bc0100000000000000000000000000000000000000040004bc0100000000000000000000000000000000000000040004bc010000000000000000000000000000000000000004000cbc010000000000000000000000000000000000000004000cbc0100000000000000000000000000000000000000040014bc0100000000000000000000000000000000000000040014bc0100000000000000000000000000000000000000040016bc0100000000000000000000000000000000000000040016bc010000000000000000000000000000000000000004001abc010000000000000000000000000000000000000004001abc0100000000000000000000000000000000000000040022bc0100000000000000000000000000000000000000040024bc0100000000000000000000000000000000000000040024bc010000000000000000000000000000000000000004002cbc010000000000000000000000000000000000000004002cbc0100000000000000000000000000000000000000040030bc0100000000000000000000000000000000000000040030bc010000000000000000000000000000000000000004003abc010000000000000000000000000000000000000004003abc0100000000000000000000000000000000000000040044bc0100000000000000000000000000473c00000000040044bc0100000000000000000000000000553c0000010001002e060100000000000200000000000000000000000000040044bc010000000000000000000000000000000000000004005abc010000000000000000000000000000000000000004005abc010000000000000000000000000000000000000004005cbc0100000000000000000000000000000000000000040060bc0100000000000000000000000000000000000000040060bc010000000000000000000000000000000000000004006ebc010000000000000000000000000000000000000004006ebc010000000000000000000000000000000000000004006ebc0100000000000000000000000000813c00000000050098c902000000000000000000000000008c3c000000000500a0c90200000000000000000000000000973c000000000500a8c90200000000000000000000000000a23c0000020004006ebc010000000000bc0100000000000000000000000004006ebc010000000000000000000000000000000000000004006ebc010000000000000000000000000000000000000004006ebc0100000000000000000000000000000000000000040070bc010000000000000000000000000000000000000004008abc01000000000000000000000000000a3d00000000040094bc0100000000000000000000000000183d0000000004009cbc0100000000000000000000000000263d000000000400a4bc01000000000000000000000000000000000000000400b4bc01000000000000000000000000000000000000000400b4bc0100000000000000000000000000343d000000000400bcbc01000000000000000000000000000000000000000400ccbc01000000000000000000000000000000000000000400ccbc01000000000000000000000000000000000000000400d0bc01000000000000000000000000000000000000000400d0bc01000000000000000000000000000000000000000400dabc01000000000000000000000000000000000000000400dabc01000000000000000000000000000000000000000400debc01000000000000000000000000000000000000000400ecbc01000000000000000000000000000000000000000400ecbc01000000000000000000000000000000000000000400f4bc01000000000000000000000000000000000000000400f4bc01000000000000000000000000000000000000000400febc01000000000000000000000000000000000000000400febc0100000000000000000000000000000000000000040006bd0100000000000000000000000000000000000000040006bd010000000000000000000000000000000000000004000cbd010000000000000000000000000000000000000004000cbd0100000000000000000000000000000000000000040010bd0100000000000000000000000000000000000000040012bd010000000000000000000000000000000000000004001ebd0100000000000000000000000000000000000000040020bd0100000000000000000000000000000000000000040026bd0100000000000000000000000000000000000000040026bd010000000000000000000000000000000000000004002ebd0100000000000000000000000000000000000000040032bd0100000000000000000000000000000000000000040032bd0100000000000000000000000000000000000000040040bd0100000000000000000000000000000000000000040046bd010000000000000000000000000000000000000004004abd010000000000000000000000000000000000000004004abd010000000000000000000000000000000000000004004ebd010000000000000000000000000000000000000004004ebd0100000000000000000000000000000000000000040054bd0100000000000000000000000000000000000000040056bd0100000000000000000000000000000000000000040056bd0100000000000000000000000000000000000000040058bd0100000000000000000000000000000000000000040058bd0100000000000000000000000000000000000000040060bd0100000000000000000000000000000000000000040060bd010000000000000000000000000000000000000004006abd010000000000000000000000000000000000000004006cbd010000000000000000000000000000000000000004006cbd010000000000000000000000000000000000000004006ebd010000000000000000000000000000000000000004006ebd0100000000000000000000000000000000000000040076bd0100000000000000000000000000000000000000040076bd0100000000000000000000000000000000000000040078bd010000000000000000000000000000000000000004007ebd010000000000000000000000000000000000000004007ebd010000000000000000000000000000000000000004008abd010000000000000000000000000000000000000004008cbd0100000000000000000000000000000000000000040090bd0100000000000000000000000000000000000000040090bd0100000000000000000000000000000000000000040094bd0100000000000000000000000000000000000000040098bd010000000000000000000000000000000000000004009ebd010000000000000000000000000000000000000004009ebd01000000000000000000000000000000000000000400aabd01000000000000000000000000000000000000000400b2bd01000000000000000000000000000000000000000400b2bd01000000000000000000000000000000000000000400b4bd01000000000000000000000000000000000000000400b6bd01000000000000000000000000000000000000000400bebd01000000000000000000000000000000000000000400bebd01000000000000000000000000000000000000000400c0bd01000000000000000000000000000000000000000400c0bd01000000000000000000000000000000000000000400c4bd01000000000000000000000000000000000000000400c4bd01000000000000000000000000000000000000000400c8bd01000000000000000000000000000000000000000400c8bd01000000000000000000000000000000000000000400dcbd01000000000000000000000000000000000000000400e2bd01000000000000000000000000000000000000000400f0bd01000000000000000000000000000000000000000400f8bd01000000000000000000000000000000000000000400f8bd01000000000000000000000000000000000000000400fcbd01000000000000000000000000000000000000000400fcbd010000000000000000000000000000000000000004000cbe0100000000000000000000000000000000000000040026be010000000000000000000000000000000000000004002abe010000000000000000000000000000000000000004002abe0100000000000000000000000000423d0000020004002abe010000000000b40000000000000000000000000004002abe010000000000000000000000000000000000000004002abe010000000000000000000000000000000000000004002abe010000000000000000000000000000000000000004002cbe010000000000000000000000000000000000000004002ebe0100000000000000000000000000000000000000040036be0100000000000000000000000000000000000000040038be0100000000000000000000000000000000000000040038be010000000000000000000000000000000000000004003cbe010000000000000000000000000000000000000004003cbe0100000000000000000000000000000000000000040044be0100000000000000000000000000000000000000040044be010000000000000000000000000000000000000004004abe010000000000000000000000000000000000000004004abe010000000000000000000000000000000000000004004ebe0100000000000000000000000000000000000000040056be010000000000000000000000000000000000000004005abe0100000000000000000000000000000000000000040066be0100000000000000000000000000000000000000040066be010000000000000000000000000000000000000004006cbe010000000000000000000000000000000000000004006cbe0100000000000000000000000000000000000000040070be0100000000000000000000000000000000000000040078be010000000000000000000000000000000000000004007ebe0100000000000000000000000000000000000000040086be010000000000000000000000000000000000000004008abe0100000000000000000000000000000000000000040096be010000000000000000000000000000000000000004009cbe01000000000000000000000000000000000000000400a4be01000000000000000000000000000000000000000400aabe01000000000000000000000000000000000000000400b2be01000000000000000000000000000000000000000400b8be01000000000000000000000000000000000000000400c0be01000000000000000000000000000000000000000400c4be01000000000000000000000000000000000000000400cebe01000000000000000000000000000000000000000400cebe01000000000000000000000000000000000000000400d8be01000000000000000000000000000000000000000400dabe01000000000000000000000000000000000000000400debe01000000000000000000000000000000000000000400debe0100000000000000000000000000753d000002000400debe01000000000038000000000000000000000000000400debe01000000000000000000000000000000000000000400debe01000000000000000000000000000000000000000400debe01000000000000000000000000000000000000000400e0be01000000000000000000000000000000000000000400e0be01000000000000000000000000000000000000000400e2be0100000000000000000000000000a63d000000000400fcbe0100000000000000000000000000b43d000001000100f8060100000000003000000000000000000000000000040010bf0100000000000000000000000000000000000000040012bf0100000000000000000000000000000000000000040016bf0100000000000000000000000000000000000000040016bf0100000000000000000000000000e03d00000200040016bf0100000000000a00000000000000000000000000040016bf0100000000000000000000000000000000000000040016bf0100000000000000000000000000000000000000040016bf0100000000000000000000000000000000000000040016bf0100000000000000000000000000000000000000040020bf0100000000000000000000000000000000000000040020bf0100000000000000000000000000363e00000200040020bf010000000000b600000000000000000000000000040020bf0100000000000000000000000000000000000000040020bf0100000000000000000000000000000000000000040020bf0100000000000000000000000000000000000000040022bf0100000000000000000000000000000000000000040022bf0100000000000000000000000000000000000000040024bf010000000000000000000000000000000000000004002ebf010000000000000000000000000000000000000004002ebf0100000000000000000000000000000000000000040030bf0100000000000000000000000000000000000000040030bf0100000000000000000000000000000000000000040034bf0100000000000000000000000000000000000000040034bf010000000000000000000000000000000000000004003cbf010000000000000000000000000000000000000004003cbf0100000000000000000000000000000000000000040042bf0100000000000000000000000000000000000000040042bf0100000000000000000000000000000000000000040046bf010000000000000000000000000000000000000004004ebf0100000000000000000000000000000000000000040052bf010000000000000000000000000000000000000004005ebf010000000000000000000000000000000000000004005ebf0100000000000000000000000000000000000000040064bf0100000000000000000000000000000000000000040064bf0100000000000000000000000000000000000000040068bf0100000000000000000000000000000000000000040070bf0100000000000000000000000000000000000000040076bf010000000000000000000000000000000000000004007ebf0100000000000000000000000000000000000000040082bf010000000000000000000000000000000000000004008ebf0100000000000000000000000000000000000000040094bf010000000000000000000000000000000000000004009cbf01000000000000000000000000000000000000000400a2bf01000000000000000000000000000000000000000400aabf01000000000000000000000000000000000000000400b0bf01000000000000000000000000000000000000000400b8bf01000000000000000000000000000000000000000400bcbf01000000000000000000000000000000000000000400c6bf01000000000000000000000000000000000000000400c6bf01000000000000000000000000000000000000000400d0bf01000000000000000000000000000000000000000400d0bf01000000000000000000000000000000000000000400d2bf01000000000000000000000000000000000000000400d6bf01000000000000000000000000000000000000000400d6bf01000000000000000000000000008e3e000002000400d6bf0100000000003a000000000000000000000000000400d6bf01000000000000000000000000000000000000000400d6bf01000000000000000000000000000000000000000400d6bf01000000000000000000000000000000000000000400d8bf01000000000000000000000000000000000000000400d8bf01000000000000000000000000000000000000000400dabf0100000000000000000000000000e43e000000000400f6bf01000000000000000000000000000000000000000400f6bf01000000000000000000000000000000000000000400f6bf010000000000000000000000000000000000000004000ac0010000000000000000000000000000000000000004000ac0010000000000000000000000000000000000000004000cc00100000000000000000000000000000000000000040010c00100000000000000000000000000000000000000040010c00100000000000000000000000000f23e00000200040010c00100000000002001000000000000000000000000040010c00100000000000000000000000000000000000000040010c00100000000000000000000000000000000000000040010c00100000000000000000000000000000000000000040012c00100000000000000000000000000000000000000040020c00100000000000000000000000000000000000000040022c00100000000000000000000000000000000000000040026c00100000000000000000000000000000000000000040026c00100000000000000000000000000000000000000040028c00100000000000000000000000000000000000000040028c00100000000000000000000000000000000000000040030c00100000000000000000000000000000000000000040034c00100000000000000000000000000000000000000040034c00100000000000000000000000000000000000000040038c00100000000000000000000000000000000000000040038c0010000000000000000000000000000000000000004003cc0010000000000000000000000000000000000000004003cc00100000000000000000000000000000000000000040040c00100000000000000000000000000000000000000040040c00100000000000000000000000000000000000000040044c00100000000000000000000000000000000000000040044c00100000000000000000000000000000000000000040046c0010000000000000000000000000000000000000004004ac001000000000000000000000000002e3f0000000004004ec001000000000000000000000000003c3f0000010001002606010000000000020000000000000000000000000004004ec00100000000000000000000000000000000000000040058c0010000000000000000000000000000000000000004005cc0010000000000000000000000000000000000000004005cc00100000000000000000000000000683f00000000040066c00100000000000000000000000000763f00000100010028060100000000000200000000000000000000000000040072c00100000000000000000000000000000000000000040072c00100000000000000000000000000000000000000040074c00100000000000000000000000000a23f0000000004007ac00100000000000000000000000000b03f0000010001002a060100000000000100000000000000000000000000040082c00100000000000000000000000000000000000000040082c0010000000000000000000000000000000000000004008cc0010000000000000000000000000000000000000004008cc0010000000000000000000000000000000000000004008ec0010000000000000000000000000000000000000004008ec00100000000000000000000000000000000000000040092c00100000000000000000000000000000000000000040092c00100000000000000000000000000000000000000040094c00100000000000000000000000000000000000000040094c001000000000000000000000000000000000000000400a0c001000000000000000000000000000000000000000400a0c001000000000000000000000000000000000000000400a4c001000000000000000000000000000000000000000400a4c001000000000000000000000000000000000000000400a6c001000000000000000000000000000000000000000400aac001000000000000000000000000000000000000000400aac001000000000000000000000000000000000000000400b2c001000000000000000000000000000000000000000400b2c001000000000000000000000000000000000000000400bcc001000000000000000000000000000000000000000400bcc001000000000000000000000000000000000000000400c0c001000000000000000000000000000000000000000400c4c001000000000000000000000000000000000000000400ccc001000000000000000000000000000000000000000400d4c001000000000000000000000000000000000000000400e8c001000000000000000000000000000000000000000400e8c001000000000000000000000000000000000000000400ecc00100000000000000000000000000dc3f000000000400ecc00100000000000000000000000000ea3f000001000100e80501000000000030000000000000000000000000000400ecc001000000000000000000000000000000000000000400f6c001000000000000000000000000000000000000000400f6c001000000000000000000000000000000000000000400fec001000000000000000000000000000000000000000400fec00100000000000000000000000000164000000000040004c10100000000000000000000000000244000000100010024060100000000000200000000000000000000000000040010c10100000000000000000000000000000000000000040010c10100000000000000000000000000000000000000040012c10100000000000000000000000000000000000000040012c10100000000000000000000000000000000000000040016c1010000000000000000000000000000000000000004001cc1010000000000000000000000000000000000000004002cc10100000000000000000000000000000000000000040030c10100000000000000000000000000000000000000040030c10100000000000000000000000000504000000200040030c10100000000000001000000000000000000000000040030c10100000000000000000000000000000000000000040030c10100000000000000000000000000000000000000040030c10100000000000000000000000000000000000000040032c10100000000000000000000000000000000000000040040c10100000000000000000000000000000000000000040042c10100000000000000000000000000000000000000040042c1010000000000000000000000000000000000000004004ac1010000000000000000000000000000000000000004004ac1010000000000000000000000000000000000000004004cc1010000000000000000000000000000000000000004004cc10100000000000000000000000000000000000000040050c10100000000000000000000000000000000000000040054c10100000000000000000000000000000000000000040054c10100000000000000000000000000000000000000040064c10100000000000000000000000000000000000000040068c1010000000000000000000000000000000000000004006cc1010000000000000000000000000000000000000004006cc10100000000000000000000000000000000000000040070c10100000000000000000000000000000000000000040070c10100000000000000000000000000000000000000040074c10100000000000000000000000000000000000000040074c10100000000000000000000000000000000000000040078c10100000000000000000000000000000000000000040078c1010000000000000000000000000000000000000004007cc1010000000000000000000000000000000000000004007cc1010000000000000000000000000000000000000004007ec10100000000000000000000000000000000000000040080c10100000000000000000000000000000000000000040080c1010000000000000000000000000089400000000004008ac10100000000000000000000000000000000000000040098c10100000000000000000000000000000000000000040098c1010000000000000000000000000000000000000004009ac101000000000000000000000000000000000000000400a4c101000000000000000000000000000000000000000400a6c101000000000000000000000000000000000000000400a6c101000000000000000000000000009740000000000400b0c10100000000000000000000000000a5400000010001002c0601000000000001000000000000000000000000000400bec101000000000000000000000000000000000000000400bec101000000000000000000000000000000000000000400c0c101000000000000000000000000000000000000000400c0c101000000000000000000000000000000000000000400c4c101000000000000000000000000000000000000000400c4c101000000000000000000000000000000000000000400c6c101000000000000000000000000000000000000000400cac101000000000000000000000000000000000000000400cac101000000000000000000000000000000000000000400d2c101000000000000000000000000000000000000000400d2c101000000000000000000000000000000000000000400dcc101000000000000000000000000000000000000000400dcc101000000000000000000000000000000000000000400e0c101000000000000000000000000000000000000000400e4c101000000000000000000000000000000000000000400ecc101000000000000000000000000000000000000000400f4c10100000000000000000000000000d14000000000040008c20100000000000000000000000000000000000000040012c20100000000000000000000000000000000000000040012c2010000000000000000000000000000000000000004001ac2010000000000000000000000000000000000000004001ac20100000000000000000000000000df4000000000040020c20100000000000000000000000000000000000000040030c20100000000000000000000000000000000000000040030c20100000000000000000000000000000000000000040030c20100000000000000000000000000000000000000040030c20100000000000000000000000000000000000000040030c20100000000000000000000000000000000000000040030c20100000000000000000000000000000000000000040032c2010000000000000000000000000000000000000004003ac2010000000000000000000000000000000000000004003cc2010000000000000000000000000000000000000004003cc20100000000000000000000000000000000000000040048c20100000000000000000000000000000000000000040048c20100000000000000000000000000000000000000040054c20100000000000000000000000000000000000000040054c20100000000000000000000000000000000000000040062c20100000000000000000000000000000000000000040062c20100000000000000000000000000000000000000040064c20100000000000000000000000000000000000000040068c2010000000000000000000000000000000000000004006ac2010000000000000000000000000000000000000004006cc2010000000000000000000000000000000000000004006cc2010000000000000000000000000000000000000004006ec2010000000000000000000000000000000000000004006ec20100000000000000000000000000000000000000040078c2010000000000000000000000000000000000000004007ac20100000000000000000000000000000000000000040082c20100000000000000000000000000000000000000040082c20100000000000000000000000000000000000000040088c20100000000000000000000000000000000000000040088c2010000000000000000000000000000000000000004008ac2010000000000000000000000000000000000000004008ac20100000000000000000000000000ed4000000000040090c20100000000000000000000000000fb400000010001002b06010000000000010000000000000000000000000004009ec2010000000000000000000000000000000000000004009ec201000000000000000000000000000000000000000400a0c201000000000000000000000000000000000000000400a0c201000000000000000000000000002741000000000400a6c201000000000000000000000000003541000001000100cc0501000000000001000000000000000000000000000400b6c201000000000000000000000000000000000000000400b6c201000000000000000000000000000000000000000400bac201000000000000000000000000000000000000000400bac201000000000000000000000000000000000000000400c4c201000000000000000000000000000000000000000400c8c201000000000000000000000000000000000000000400c8c201000000000000000000000000000000000000000400c8c201000000000000000000000000000000000000000400c8c201000000000000000000000000000000000000000400c8c201000000000000000000000000000000000000000400cac201000000000000000000000000000000000000000400cac201000000000000000000000000000000000000000400ccc201000000000000000000000000000000000000000400d6c201000000000000000000000000000000000000000400d6c201000000000000000000000000006141000002000400d6c201000000000072000000000000000000000000000400d6c201000000000000000000000000000000000000000400d6c201000000000000000000000000000000000000000400d6c201000000000000000000000000000000000000000400d8c201000000000000000000000000000000000000000400dac201000000000000000000000000000000000000000400dcc201000000000000000000000000000000000000000400dcc201000000000000000000000000000000000000000400e4c201000000000000000000000000000000000000000400e4c201000000000000000000000000000000000000000400f0c201000000000000000000000000000000000000000400f0c201000000000000000000000000000000000000000400f2c201000000000000000000000000000000000000000400f2c201000000000000000000000000000000000000000400f6c201000000000000000000000000000000000000000400f6c201000000000000000000000000000000000000000400fec201000000000000000000000000000000000000000400fec20100000000000000000000000000000000000000040006c30100000000000000000000000000000000000000040006c3010000000000000000000000000000000000000004000ac3010000000000000000000000000000000000000004000ac30100000000000000000000000000000000000000040014c30100000000000000000000000000000000000000040014c3010000000000000000000000000000000000000004001ec30100000000000000000000000000c0410000000004001ec3010000000000000000000000000000000000000004001ec30100000000000000000000000000000000000000040034c30100000000000000000000000000000000000000040034c30100000000000000000000000000000000000000040036c3010000000000000000000000000000000000000004003ac3010000000000000000000000000000000000000004003ac30100000000000000000000000000000000000000040048c30100000000000000000000000000000000000000040048c30100000000000000000000000000000000000000040048c30100000000000000000000000000ce4100000200040048c30100000000007200000000000000000000000000040048c30100000000000000000000000000000000000000040048c30100000000000000000000000000000000000000040048c3010000000000000000000000000000000000000004004ac3010000000000000000000000000000000000000004004cc3010000000000000000000000000000000000000004004ec3010000000000000000000000000000000000000004004ec30100000000000000000000000000000000000000040056c30100000000000000000000000000000000000000040056c30100000000000000000000000000000000000000040062c30100000000000000000000000000000000000000040062c30100000000000000000000000000000000000000040064c30100000000000000000000000000000000000000040064c30100000000000000000000000000000000000000040068c30100000000000000000000000000000000000000040068c30100000000000000000000000000000000000000040070c30100000000000000000000000000000000000000040070c30100000000000000000000000000000000000000040078c30100000000000000000000000000000000000000040078c3010000000000000000000000000000000000000004007cc3010000000000000000000000000000000000000004007cc30100000000000000000000000000000000000000040086c30100000000000000000000000000000000000000040086c30100000000000000000000000000000000000000040090c301000000000000000000000000002d4200000000040090c30100000000000000000000000000000000000000040090c301000000000000000000000000000000000000000400a6c301000000000000000000000000000000000000000400a6c301000000000000000000000000000000000000000400a8c301000000000000000000000000000000000000000400acc301000000000000000000000000000000000000000400acc301000000000000000000000000000000000000000400bac301000000000000000000000000000000000000000400bac301000000000000000000000000000000000000000400bac301000000000000000000000000003b42000002000400bac301000000000016000000000000000000000000000400bac301000000000000000000000000000000000000000400bac301000000000000000000000000008342000000000400bac301000000000000000000000000000000000000000400bac301000000000000000000000000009142000001000100280701000000000002000000000000000000000000000400bac301000000000000000000000000000000000000000400d0c301000000000000000000000000000000000000000400d0c301000000000000000000000000000000000000000400d0c30100000000000000000000000000bd42000002000400d0c3010000000000a2000000000000000000000000000400d0c301000000000000000000000000000000000000000400d0c301000000000000000000000000000000000000000400d0c301000000000000000000000000000000000000000400d2c301000000000000000000000000000000000000000400d8c301000000000000000000000000000000000000000400dac301000000000000000000000000000000000000000400dac301000000000000000000000000000000000000000400dcc301000000000000000000000000000000000000000400dcc301000000000000000000000000000000000000000400dec301000000000000000000000000000000000000000400dec301000000000000000000000000001e43000000000400e2c301000000000000000000000000002c43000001000100500701000000000011000000000000000000000000000400eec301000000000000000000000000000000000000000400eec301000000000000000000000000000000000000000400fac301000000000000000000000000005843000000000400fac301000000000000000000000000006643000001000100300701000000000020000000000000000000000000000400fac3010000000000000000000000000000000000000004000ec4010000000000000000000000000000000000000004000ec40100000000000000000000000000000000000000040010c40100000000000000000000000000000000000000040014c40100000000000000000000000000000000000000040016c40100000000000000000000000000000000000000040018c40100000000000000000000000000000000000000040018c4010000000000000000000000000000000000000004001ac4010000000000000000000000000000000000000004001ac40100000000000000000000000000000000000000040024c40100000000000000000000000000000000000000040026c4010000000000000000000000000000000000000004002ec4010000000000000000000000000000000000000004002ec40100000000000000000000000000000000000000040034c40100000000000000000000000000000000000000040034c40100000000000000000000000000000000000000040036c40100000000000000000000000000000000000000040036c4010000000000000000000000000092430000000004003cc4010000000000000000000000000000000000000004004ac4010000000000000000000000000000000000000004004ac4010000000000000000000000000000000000000004004cc4010000000000000000000000000000000000000004004cc40100000000000000000000000000a04300000000040052c40100000000000000000000000000000000000000040062c40100000000000000000000000000000000000000040062c40100000000000000000000000000000000000000040066c40100000000000000000000000000000000000000040066c4010000000000000000000000000000000000000004006ec40100000000000000000000000000000000000000040072c40100000000000000000000000000000000000000040072c40100000000000000000000000000ae4300000200040072c40100000000007000000000000000000000000000040072c40100000000000000000000000000000000000000040072c40100000000000000000000000000000000000000040072c40100000000000000000000000000000000000000040074c40100000000000000000000000000000000000000040076c40100000000000000000000000000000000000000040078c40100000000000000000000000000000000000000040078c40100000000000000000000000000000000000000040080c40100000000000000000000000000000000000000040080c40100000000000000000000000000000000000000040088c40100000000000000000000000000000000000000040088c4010000000000000000000000000000000000000004008ac4010000000000000000000000000000000000000004008ac4010000000000000000000000000000000000000004008ec4010000000000000000000000000000000000000004008ec40100000000000000000000000000000000000000040096c40100000000000000000000000000000000000000040098c40100000000000000000000000000000000000000040098c401000000000000000000000000000000000000000400a0c401000000000000000000000000000000000000000400a0c401000000000000000000000000000000000000000400a4c401000000000000000000000000000000000000000400a4c401000000000000000000000000000000000000000400aec401000000000000000000000000000000000000000400aec401000000000000000000000000000000000000000400b8c401000000000000000000000000000e44000000000400b8c401000000000000000000000000000000000000000400b8c401000000000000000000000000000000000000000400cec401000000000000000000000000000000000000000400cec401000000000000000000000000000000000000000400d0c401000000000000000000000000000000000000000400d4c401000000000000000000000000000000000000000400d4c401000000000000000000000000000000000000000400e2c401000000000000000000000000000000000000000400e2c401000000000000000000000000000000000000000400e2c401000000000000000000000000000000000000000400e2c401000000000000000000000000000000000000000400e4c401000000000000000000000000000000000000000400eec401000000000000000000000000001c4400000200040034c50100000000007e00000000000000000000000000040034c50100000000000000000000000000000000000000040034c50100000000000000000000000000000000000000040036c5010000000000000000000000000000000000000004003cc501000000000000000000000000000000000000000400b2c501000000000000000000000000000000000000000400b2c501000000000000000000000000000000000000000400b4c501000000000000000000000000000000000000000400bcc50100000000000000000000000000000000000000040014c60100000000000000000000000000764400000200040014c60100000000003600000000000000000000000000040014c6010000000000000000000000000000000000000004004ac60100000000000000000000000000be440000020004004ac6010000000000300000000000000000000000000004004ac6010000000000000000000000000000000000000004007ac6010000000000000000000000000000000000000004007ac6010000000000000000000000000000000000000004007cc60100000000000000000000000000000000000000040080c601000000000000000000000000000000000000000400c8c601000000000000000000000000000645000002000400c8c601000000000086000000000000000000000000000400c8c601000000000000000000000000000000000000000400cac601000000000000000000000000000000000000000400d6c601000000000000000000000000006545000000000400e4c601000000000000000000000000007345000001000100e60501000000000001000000000000009f45000000000400fec60100000000000000000000000000ad450000000004002ec70100000000000000000000000000bb450000010001002d06010000000000010000000000000000000000000004004ec70100000000000000000000000000e7450000020004004ec7010000000000680000000000000000000000000004004ec70100000000000000000000000000000000000000040050c7010000000000000000000000000000000000000004005ac701000000000000000000000000002846000002000400b6c70100000000007e000000000000000000000000000400b6c701000000000000000000000000000000000000000400b6c701000000000000000000000000000000000000000400b8c701000000000000000000000000000000000000000400bec70100000000000000000000000000824600000200040034c80100000000005200000000000000000000000000040034c80100000000000000000000000000000000000000040034c80100000000000000000000000000000000000000040036c8010000000000000000000000000000000000000004003cc80100000000000000000000000000000000000000040086c80100000000000000000000000000000000000000040086c80100000000000000000000000000000000000000040088c8010000000000000000000000000000000000000004008cc801000000000000000000000000000000000000000400dcc80100000000000000000000000000b546000002000400dcc801000000000082010000000000000000000000000400dcc801000000000000000000000000000000000000000400dec801000000000000000000000000000000000000000400ecc80100000000000000000000000000e646000000000400bec90100000000000000000000000000f44600000100010000080100000000001c00000000000000fe46000000000400c8c901000000000000000000000000000c47000000000400d2c901000000000000000000000000001a47000000000400e6c901000000000000000000000000002847000000000400eec901000000000000000000000000003647000001000100880701000000000020000000000000006047000000000400fcc901000000000000000000000000006e4700000100010066080100000000002f0000000000000099470000000004000aca0100000000000000000000000000a74700000100010095080100000000003200000000000000d24700000000040024ca0100000000000000000000000000e0470000000004002cca0100000000000000000000000000ee47000001000100e0070100000000002000000000000000184800000000040046ca010000000000000000000000000026480000010001001c080100000000001c00000000000000514800000000040050ca01000000000000000000000000005f4800000100010038080100000000002e0000000000000000000000000004005eca01000000000000000000000000008a480000020004005eca010000000000280000000000000000000000000004005eca0100000000000000000000000000e54800000000040064ca0100000000000000000000000000f348000001000100d00d01000000000050000000000000005d490000000004006eca01000000000000000000000000006b49000001000100200e0100000000005000000000000000000000000000040086ca0100000000000000000000000000000000000000040086ca0100000000000000000000000000000000000000040088ca0100000000000000000000000000d949000000000400a8ca0100000000000000000000000000e749000000000400b4ca0100000000000000000000000000f549000001000100a80701000000000018000000000000001f4a000000000400bcca01000000000000000000000000002d4a000001000100c0070100000000002000000000000000574a000000000400d2ca0100000000000000000000000000654a000001000100c70801000000000026000000000000000000000000000400e8ca0100000000000000000000000000904a000002000400e8ca01000000000068000000000000000000000000000400e8ca01000000000000000000000000000000000000000400eaca01000000000000000000000000000000000000000400eeca0100000000000000000000000000cf4a0000000004001acb0100000000000000000000000000dd4a00000000040022cb0100000000000000000000000000eb4a0000000004003ccb0100000000000000000000000000f94a000001000100ed080100000000000d00000000000000000000000000040050cb0100000000000000000000000000000000000000040050cb0100000000000000000000000000000000000000040052cb0100000000000000000000000000000000000000040054cb0100000000000000000000000000244b0000000004006ccb0100000000000000000000000000324b000001000100fa080100000000000e00000000000000000000000000040080cb0100000000000000000000000000000000000000040080cb0100000000000000000000000000000000000000040082cb0100000000000000000000000000000000000000040094cb01000000000000000000000000005d4b00000000040010cc01000000000000000000000000006b4b0000000004009ecc0100000000000000000000000000794b000000000400a8cc0100000000000000000000000000874b000000000400b2cc0100000000000000000000000000954b000000000400bccc0100000000000000000000000000a34b000000000400c6cc0100000000000000000000000000b14b000000000400d0cc01000000000000000000000000000000000000000400e6cc01000000000000000000000000000000000000000400e6cc01000000000000000000000000000000000000000400e8cc01000000000000000000000000000000000000000400eccc0100000000000000000000000000bf4b00000000040034cd010000000000000000000000000000000000000004004acd010000000000000000000000000000000000000004004acd010000000000000000000000000000000000000004004ccd0100000000000000000000000000000000000000040052cd0100000000000000000000000000cd4b0000000004008ccd0100000000000000000000000000db4b00000000040094cd0100000000000000000000000000e94b000000000400aecd0100000000000000000000000000f74b00000100010008090100000000000e000000000000000000000000000400c2cd01000000000000000000000000000000000000000400c2cd01000000000000000000000000000000000000000400c4cd01000000000000000000000000000000000000000400cacd0100000000000000000000000000224c0000000004000ace0100000000000000000000000000304c00000000040012ce01000000000000000000000000003e4c0000000004002cce01000000000000000000000000004c4c00000100010024090100000000000d00000000000000000000000000040040ce0100000000000000000000000000000000000000040040ce0100000000000000000000000000000000000000040042ce010000000000000000000000000000000000000004004ace0100000000000000000000000000774c000000000400acce0100000000000000000000000000854c000000000400b4ce0100000000000000000000000000934c000000000400cece0100000000000000000000000000a14c000001000100310901000000000012000000000000000000000000000400e2ce0100000000000000000000000000cc4c000002000400e2ce0100000000007a000000000000000000000000000400e2ce01000000000000000000000000000000000000000400e4ce01000000000000000000000000000000000000000400eace0100000000000000000000000000304d0000000004003acf010000000000000000000000000000000000000004005ccf010000000000000000000000000000000000000004005ccf010000000000000000000000000000000000000004005ecf010000000000000000000000000000000000000004006acf01000000000000000000000000003e4d000000000400c4cf01000000000000000000000000004c4d00000100010048090100000000002000000000000000000000000000040016d00100000000000000000000000000774d00000200040016d00100000000001000000000000000000000000000040016d00100000000000000000000000000000000000000040026d00100000000000000000000000000c84d00000200040026d00100000000008c00000000000000000000000000040026d00100000000000000000000000000000000000000040028d00100000000000000000000000000000000000000040030d001000000000000000000000000000000000000000400b2d001000000000000000000000000000b4e000002000400b2d00100000000004a000000000000000000000000000400b2d001000000000000000000000000000000000000000400fcd001000000000000000000000000006f4e000002000400fcd001000000000072000000000000000000000000000400fcd001000000000000000000000000000000000000000400fed00100000000000000000000000000000000000000040006d10100000000000000000000000000f04e00000000040050d10100000000000000000000000000fe4e000001000100100a0100000000001c0000000000000000000000000004006ed1010000000000000000000000000000000000000004006ed10100000000000000000000000000084f0000000004000ed20100000000000000000000000000164f00000000040024d2010000000000000000000000000000000000000004002ed20100000000000000000000000000244f0000020004002ed2010000000000280000000000000000000000000004002ed20100000000000000000000000000000000000000040030d20100000000000000000000000000000000000000040032d20100000000000000000000000000000000000000040056d20100000000000000000000000000694f00000200040056d20100000000002800000000000000000000000000040056d20100000000000000000000000000000000000000040058d2010000000000000000000000000000000000000004005ad2010000000000000000000000000000000000000004007ed20100000000000000000000000000ae4f0000020004007ed2010000000000140100000000000000000000000004007ed20100000000000000000000000000000000000000040080d20100000000000000000000000000000000000000040098d20100000000000000000000000000000000000000040092d30100000000000000000000000000c95000000200040092d30100000000006c00000000000000000000000000040092d301000000000000000000000000000000000000000400fed301000000000000000000000000006e51000002000400fed30100000000007e030000000000000000000000000400fed30100000000000000000000000000000000000000040000d4010000000000000000000000000000000000000004001ad40100000000000000000000000000bc5200000200040082da010000000000e8020000000000002c530000020004007cd7010000000000060300000000000093530000020004006add010000000000d002000000000000f9530000020004003ae0010000000000ae0200000000000000000000000004007cd7010000000000000000000000000000000000000004007cd7010000000000000000000000000000000000000004007ed70100000000000000000000000000000000000000040098d7010000000000000000000000000057540000000004003eda010000000000000000000000000065540000010001009e0b0100000000001b0000000000000090540000000004004ada01000000000000000000000000009e5400000000040058da0100000000000000000000000000ac5400000000040062da0100000000000000000000000000ba540000000004006cda0100000000000000000000000000000000000000040082da0100000000000000000000000000000000000000040082da0100000000000000000000000000000000000000040084da010000000000000000000000000000000000000004009eda0100000000000000000000000000c85400000000040046dd0100000000000000000000000000d65400000000040054dd010000000000000000000000000000000000000004006add010000000000000000000000000000000000000004006add010000000000000000000000000000000000000004006cdd0100000000000000000000000000000000000000040086dd0100000000000000000000000000e454000000000400f2df0100000000000000000000000000f254000000000400fedf010000000000000000000000000000550000000004000ce001000000000000000000000000000e550000000004001ae001000000000000000000000000001c5500000000040024e0010000000000000000000000000000000000000004003ae0010000000000000000000000000000000000000004003ae0010000000000000000000000000000000000000004003ce00100000000000000000000000000000000000000040056e001000000000000000000000000002a55000000000400d2e201000000000000000000000000000000000000000400e8e201000000000000000000000000003855000002000400e8e201000000000028000000000000000000000000000400e8e201000000000000000000000000000000000000000400eae201000000000000000000000000000000000000000400ece20100000000000000000000000000000000000000040010e301000000000000000000000000007d5500000200040010e30100000000002800000000000000000000000000040010e30100000000000000000000000000000000000000040012e30100000000000000000000000000000000000000040014e30100000000000000000000000000000000000000040038e30100000000000000000000000000c25500000200040038e30100000000002801000000000000000000000000040038e3010000000000000000000000000000000000000004003ae30100000000000000000000000000000000000000040050e30100000000000000000000000000000000000000040060e40100000000000000000000000000dd5600000200040060e40100000000006800000000000000000000000000040060e40100000000000000000000000000000000000000040062e40100000000000000000000000000000000000000040070e401000000000000000000000000000000000000000400c8e401000000000000000000000000008257000002000400c8e401000000000004030000000000000000000000000400c8e401000000000000000000000000000000000000000400cce40100000000000000000000000000000000000000040000e50100000000000000000000000000d058000002000400cce701000000000066000000000000009859000002000400f8ea0100000000004602000000000000085a00000200040032e8010000000000c6020000000000006f5a0000020004003eed0100000000008e02000000000000d55a000002000400ccef01000000000002020000000000000000000000000400cce701000000000000000000000000000000000000000400cce70100000000000000000000000000000000000000040032e80100000000000000000000000000000000000000040032e80100000000000000000000000000000000000000040036e8010000000000000000000000000000000000000004006ae80100000000000000000000000000335b000000000400b4ea0100000000000000000000000000415b000000000400c0ea01000000000000000000000000004f5b000000000400ceea01000000000000000000000000005d5b000000000400d8ea01000000000000000000000000006b5b000000000400e2ea01000000000000000000000000000000000000000400f8ea01000000000000000000000000000000000000000400f8ea01000000000000000000000000000000000000000400faea0100000000000000000000000000000000000000040014eb0100000000000000000000000000795b0000000004001aed0100000000000000000000000000875b00000000040028ed010000000000000000000000000000000000000004003eed010000000000000000000000000000000000000004003eed0100000000000000000000000000000000000000040042ed0100000000000000000000000000000000000000040076ed0100000000000000000000000000955b00000000040084ef0100000000000000000000000000a35b00000000040090ef0100000000000000000000000000b15b0000000004009eef0100000000000000000000000000bf5b000000000400acef0100000000000000000000000000cd5b000000000400b6ef01000000000000000000000000000000000000000400ccef01000000000000000000000000000000000000000400ccef01000000000000000000000000000000000000000400ceef01000000000000000000000000000000000000000400e8ef0100000000000000000000000000db5b000000000400b8f101000000000000000000000000000000000000000400cef10100000000000000000000000000e95b000002000400cef101000000000036290000000000000000000000000400cef101000000000000000000000000000000000000000400d2f101000000000000000000000000000000000000000400fcf10100000000000000000000000000195c000002000400a82002000000000006040000000000005c5c000002000400962e0200000000005001000000000000945c000002000400e62f0200000000000c03000000000000d45c000002000400ae24020000000000e8090000000000000000000000000400041b0200000000000000000000000000055d000000000500b0c90200000000000000000000000000105d000002000400041b0200000000008e000000000000000000000000000400041b02000000000000000000000000000000000000000400061b020000000000000000000000000000000000000004000c1b02000000000000000000000000005d5d000000000400261b02000000000000000000000000000000000000000400921b02000000000000000000000000006b5d000002000400921b020000000000cc010000000000000000000000000400921b02000000000000000000000000000000000000000400961b02000000000000000000000000000000000000000400ae1b0200000000000000000000000000a35d000000000400c81b0200000000000000000000000000b15d000002000400ba360200000000006a00000000000000df5d0000020004005e1d020000000000f600000000000000225e000000000400b81c0200000000000000000000000000305e000000000400dc1c02000000000000000000000000003e5e000002000400541e020000000000540200000000000000000000000004005e1d020000000000000000000000000000000000000004005e1d02000000000000000000000000000000000000000400621d02000000000000000000000000000000000000000400761d02000000000000000000000000000000000000000400541e02000000000000000000000000000000000000000400541e02000000000000000000000000000000000000000400581e02000000000000000000000000000000000000000400701e02000000000000000000000000000000000000000400a82002000000000000000000000000000000000000000400a82002000000000000000000000000000000000000000400aa2002000000000000000000000000000000000000000400c0200200000000000000000000000000815e000000000400982402000000000000000000000000008f5e000001000100300a0100000000002e000000000000000000000000000400ae2402000000000000000000000000000000000000000400ae2402000000000000000000000000000000000000000400b02402000000000000000000000000000000000000000400c82402000000000000000000000000000000000000000400962e0200000000000000000000000000ba5e000000000500b8c90200000000000000000000000000c55e000000000500c0c90200000000000000000000000000d05e000000000500c8c90200000000000000000000000000db5e000000000500d0c902000000000000000000000000000000000000000400962e02000000000000000000000000000000000000000400982e02000000000000000000000000000000000000000400aa2e0200000000000000000000000000e65e000000000400d62e0200000000000000000000000000f45e000000000400de2e0200000000000000000000000000025f000000000400f82e0200000000000000000000000000105f000000000400002f02000000000000000000000000001e5f000000000400d22f02000000000000000000000000000000000000000400e62f02000000000000000000000000000000000000000400e62f02000000000000000000000000000000000000000400e82f02000000000000000000000000000000000000000400023002000000000000000000000000002c5f000002000400f232020000000000c8030000000000000000000000000400f23202000000000000000000000000000000000000000400f23202000000000000000000000000000000000000000400f43202000000000000000000000000000000000000000400043302000000000000000000000000000000000000000400ba3602000000000000000000000000000000000000000400ba3602000000000000000000000000000000000000000400bc3602000000000000000000000000000000000000000400c4360200000000000000000000000000705f000000000400ec3602000000000000000000000000000000000000000400243702000000000000000000000000007e5f000000000500d8c90200000000000000000000000000895f00000200040024370200000000008e0000000000000000000000000004002437020000000000000000000000000000000000000004002637020000000000000000000000000000000000000004002c370200000000000000000000000000d65f000000000400463702000000000000000000000000000000000000000400b2370200000000000000000000000000e45f000002000400b23702000000000072000000000000000000000000000400b23702000000000000000000000000000000000000000400b43702000000000000000000000000000000000000000400bc3702000000000000000000000000006560000000000400103802000000000000000000000000000000000000000400243802000000000000000000000000000000000000000400243802000000000000000000000000007360000000000400263802000000000000000000000000008160000000000100880101000000000000000000000000008c6000000000040036380200000000000000000000000000966000000000040038380200000000000000000000000000a0600000000004003a380200000000000000000000000000aa600000000004003e380200000000000000000000000000b4600000000004004238020000000000000000000000000000000000000004004c38020000000000000000000000000000000000000004004c38020000000000000000000000000000000000000004006838020000000000000000000000000000000000000004006838020000000000000000000000000000000000000004006c380200000000000000000000000000000000000000040084380200000000000000000000000000be60000000000400ba380200000000000000000000000000000000000000040042390200000000000000000000000000000000000000040042390200000000000000000000000000000000000000040044390200000000000000000000000000000000000000040050390200000000000000000000000000cc600000020004006c3b02000000000032000000000000003e610000000004004c3b02000000000000000000000000004c61000000000400543b02000000000000000000000000005a61000001000100900a010000000000200000000000000000000000000004006c3b020000000000000000000000000000000000000004006c3b020000000000000000000000000000000000000004006e3b02000000000000000000000000000000000000000400723b020000000000000000000000000000000000000004009e3b020000000000000000000000000000000000000004009e3b02000000000000000000000000000000000000000400a03b02000000000000000000000000000000000000000400b63b02000000000000000000000000008561000000000400743e02000000000000000000000000009361000000000400883e0200000000000000000000000000a161000001000100500d0100000000002b00000000000000cd61000000000400963e0200000000000000000000000000db610000000004009e3e02000000000000000000000000000000000000000400b63e02000000000000000000000000000000000000000400b63e02000000000000000000000000000000000000000400b83e02000000000000000000000000000000000000000400d23e0200000000000000000000000000e96100000000040000420200000000000000000000000000f7610000000004001442020000000000000000000000000005620000000004001c4202000000000000000000000000001362000001000100b00a01000000000020000000000000003e62000000000400344202000000000000000000000000004c620000010001007b0d010000000000290000000000000000000000000004004242020000000000000000000000000000000000000004004242020000000000000000000000000000000000000004004442020000000000000000000000000000000000000004005e4202000000000000000000000000007862000000000400904502000000000000000000000000008662000000000400a44502000000000000000000000000009462000000000400ac450200000000000000000000000000a262000000000400c4450200000000000000000000000000b062000001000100a40d0100000000002c000000000000000000000000000400d24502000000000000000000000000000000000000000400d24502000000000000000000000000000000000000000400d44502000000000000000000000000000000000000000400ee450200000000000000000000000000dc620000000004009e490200000000000000000000000000ea62000000000400b2490200000000000000000000000000f862000000000400ba4902000000000000000000000000000663000000000400ca4902000000000000000000000000001463000000000400d24902000000000000000000000000002263000000000400e24902000000000000000000000000003063000000000400ea4902000000000000000000000000003e63000000000400f44902000000000000000000000000004c63000000000400fc4902000000000000000000000000000000000000000400204a02000000000000000000000000000000000000000400204a02000000000000000000000000000000000000000400224a020000000000000000000000000000000000000004002e4a02000000000000000000000000005a63000000000400804b02000000000000000000000000000000000000000400a64b02000000000000000000000000006863000002000400a64b02000000000056020000000000000000000000000400a64b02000000000000000000000000000000000000000400a84b02000000000000000000000000000000000000000400c24b0200000000000000000000000000a863000000000400c84d0200000000000000000000000000b663000000000400dc4d0200000000000000000000000000c463000000000400e44d02000000000000000000000000000000000000000400fc4d02000000000000000000000000000000000000000400fc4d02000000000000000000000000000000000000000400fe4d02000000000000000000000000000000000000000400064e0200000000000000000000000000d263000000000400744e0200000000000000000000000000e0630000000004007c4e02000000000000000000000000000000000000000400964e02000000000000000000000000000000000000000400964e02000000000000000000000000000000000000000400984e020000000000000000000000000000000000000004009e4e0200000000000000000000000000ee63000000000400964f0200000000000000000000000000fc630000000004009e4f02000000000000000000000000000a64000000000400a84f02000000000000000000000000001864000000000400b04f02000000000000000000000000002664000000000400c04f02000000000000000000000000003464000000000400c84f02000000000000000000000000004264000000000400d84f02000000000000000000000000005064000000000400e04f02000000000000000000000000005e64000000000400fa4f02000000000000000000000000006c6400000100010016090100000000000e0000000000000000000000000004000e50020000000000000000000000000000000000000004000e50020000000000000000000000000000000000000004001050020000000000000000000000000000000000000004002a500200000000000000000000000000976400000000040020520200000000000000000000000000a56400000000040034520200000000000000000000000000b3640000000004003c520200000000000000000000000000c1640000000004005452020000000000000000000000000000000000000004006252020000000000000000000000000000000000000004006252020000000000000000000000000000000000000004006652020000000000000000000000000000000000000004009a520200000000000000000000000000cf64000000000400c8580200000000000000000000000000dd640000000004008a590200000000000000000000000000eb6400000100010080020100000000001c00000000000000f164000000000400b4590200000000000000000000000000ff64000000000400bc5902000000000000000000000000000d65000001000100d00a01000000000020000000000000000000000000000400d45902000000000000000000000000000000000000000400d45902000000000000000000000000000000000000000400d85902000000000000000000000000000000000000000400e45902000000000000000000000000000000000000000400485a02000000000000000000000000000000000000000400485a020000000000000000000000000000000000000004004c5a02000000000000000000000000000000000000000400805a02000000000000000000000000000000000000000400805a02000000000000000000000000000000000000000400825a02000000000000000000000000003865000000000400dc5b02000000000000000000000000004665000000000400967502000000000000000000000000005465000000000400b87502000000000000000000000000006265000000000400228802000000000000000000000000007065000000000100b00101000000000000000000000000007b650000000004000093020000000000000000000000000087650000000004005688020000000000000000000000000093650000000004002a8a02000000000000000000000000009f650000000004008e8c0200000000000000000000000000ab650000000004004a8e0200000000000000000000000000b7650000000004009a8e0200000000000000000000000000c36500000000040018930200000000000000000000000000d1650000000004002a930200000000000000000000000000df6500000000040038930200000000000000000000000000ed6500000000040046930200000000000000000000000000fb650000000004005093020000000000000000000000000009660000000004005a93020000000000000000000000000017660000000004006493020000000000000000000000000025660000000004007e93020000000000000000000000000033660000000004009493020000000000000000000000000041660000000004009e9302000000000000000000000000004f66000000000400ac9302000000000000000000000000005d66000000000400c09302000000000000000000000000006b66000000000400ca9302000000000000000000000000007966000000000400d49302000000000000000000000000008766000000000400de9302000000000000000000000000009566000000000400e8930200000000000000000000000000a366000000000400f2930200000000000000000000000000b16600000000040006940200000000000000000000000000bf6600000000040010940200000000000000000000000000cd660000000004001a940200000000000000000000000000db6600000000040024940200000000000000000000000000e9660000000004002e940200000000000000000000000000f7660000000004003894020000000000000000000000000005670000000004005a94020000000000000000000000000013670000000004006494020000000000000000000000000021670000000004006e9402000000000000000000000000002f670000000004007e9402000000000000000000000000003d67000000000400889402000000000000000000000000000000000000000400929402000000000000000000000000004b67000001000800a0ca02000000000000100800000000007a67000001000800a0da0a00000000000010000000000000af67000001000100dc030100000000002300000000000000da6700000100010010040100000000003300000000000000056800000100010068090100000000000a00000000000000306800000100010072090100000000000a000000000000005b680000010001007c090100000000000b00000000000000866800000100010087090100000000000600000000000000b1680000010001008d090100000000000600000000000000dc680000010001009309010000000000090000000000000007690000010001009c0901000000000006000000000000000000000000000a00000000000000000000000000000000000000000000000d00752b00000000000000000000000000000000000000000d00604600000000000000000000000000003269000000001100000000000000000000000000000000000000000000000d002b1300000000000000000000000000000000000000000c00701100000000000000000000000000000000000000000d00742f00000000000000000000000000000000000000000d00000000000000000000000000000000000000000000000d007c4f00000000000000000000000000000000000000000d00643800000000000000000000000000000000000000000d00953f00000000000000000000000000000000000000000d00190f00000000000000000000000000000000000000000a00740000000000000000000000000000000000000000000d005a1700000000000000000000000000004669000000001100880000000000000000000000000000000000000000000c00a01100000000000000000000000000000000000000000d003b1a00000000000000000000000000000000000000000d00840500000000000000000000000000000000000000000d002f0d00000000000000000000000000000000000000000d00901700000000000000000000000000000000000000000d00dc3500000000000000000000000000000000000000000d00dd0c00000000000000000000000000000000000000000d00ab3f00000000000000000000000000000000000000000d00973300000000000000000000000000000000000000000d00e63800000000000000000000000000000000000000000d00182500000000000000000000000000000000000000000d009a2a00000000000000000000000000000000000000000d006c2300000000000000000000000000000000000000000d00eb2c00000000000000000000000000000000000000000d00d14900000000000000000000000000000000000000000d00ba3b00000000000000000000000000000000000000000d006f3a00000000000000000000000000000000000000000d00770c00000000000000000000000000000000000000000d00f90300000000000000000000000000000000000000000d005f0d00000000000000000000000000000000000000000d00ae4200000000000000000000000000000000000000000d00b03300000000000000000000000000000000000000000d008d1800000000000000000000000000000000000000000d00ff0b00000000000000000000000000000000000000000d00d53700000000000000000000000000000000000000000d00a60000000000000000000000000000000000000000000d00794a00000000000000000000000000000000000000000d00fd1300000000000000000000000000000000000000000d00574400000000000000000000000000000000000000000d00244900000000000000000000000000000000000000000d00900500000000000000000000000000000000000000000d00b80800000000000000000000000000000000000000000d00cc0000000000000000000000000000000000000000000d000b2a00000000000000000000000000000000000000000d00933300000000000000000000000000000000000000000d005b1300000000000000000000000000000000000000000d00903400000000000000000000000000000000000000000d00fd4b00000000000000000000000000000000000000000d00542900000000000000000000000000000000000000000d007b4100000000000000000000000000000000000000000d00361400000000000000000000000000000000000000000d00c84900000000000000000000000000000000000000000d008f3e00000000000000000000000000000000000000000d00544c00000000000000000000000000000000000000000d004f3100000000000000000000000000000000000000000d00fc1600000000000000000000000000000000000000000d00763800000000000000000000000000000000000000000c00000000000000000000000000000000000000000000000c00400000000000000000000000000000000000000000000c00700000000000000000000000000000000000000000000c00a00000000000000000000000000000000000000000000d00550c00000000000000000000000000000000000000000d00472d00000000000000000000000000000000000000000d00c03e00000000000000000000000000000000000000000d00441b00000000000000000000000000000000000000000d00f20400000000000000000000000000000000000000000d00c11600000000000000000000000000000000000000000d00b41000000000000000000000000000000000000000000d00aa3000000000000000000000000000000000000000000d004e2b00000000000000000000000000000000000000000d002a2b00000000000000000000000000000000000000000d00011500000000000000000000000000000000000000000d00581d00000000000000000000000000000000000000000d008b4700000000000000000000000000000000000000000d00c54a00000000000000000000000000000000000000000d001d3c00000000000000000000000000000000000000000d00761500000000000000000000000000000000000000000d00ef3000000000000000000000000000000000000000000c00200900000000000000000000000000000000000000000c00500900000000000000000000000000000000000000000c00800900000000000000000000000000000000000000000c00b00900000000000000000000000000000000000000000c00e00900000000000000000000000000000000000000000d00c60700000000000000000000000000000000000000000d00733500000000000000000000000000000000000000000d000f0f00000000000000000000000000000000000000000d00f52800000000000000000000000000000000000000000c00100e00000000000000000000000000000000000000000c00400e00000000000000000000000000000000000000000c00700e00000000000000000000000000000000000000000c00a00e00000000000000000000000000000000000000000c00d00e00000000000000000000000000000000000000000d004b4800000000000000000000000000000000000000000d00af4800000000000000000000000000000000000000000c00000f00000000000000000000000000000000000000000c00300f00000000000000000000000000000000000000000c00600f00000000000000000000000000000000000000000c00900f00000000000000000000000000000000000000000c00c00f00000000000000000000000000000000000000000d00210800000000000000000000000000000000000000000d001f0300000000000000000000000000000000000000000c00801000000000000000000000000000000000000000000c00b01000000000000000000000000000000000000000000c00e01000000000000000000000000000000000000000000c00101100000000000000000000000000000000000000000c00401100000000000000000000000000000000000000000d00d74d00000000000000000000000000000000000000000d00e90a00000000000000000000000000000000000000000d001e0b00000000000000000000000000000000000000000d007f0300000000000000000000000000000000000000000d00533100000000000000000000000000000000000000000d00c94c00000000000000000000000000000000000000000d00434400000000000000000000000000000000000000000d006b0d00000000000000000000000000000000000000000d00880500000000000000000000000000000000000000000d00890200000000000000000000000000000000000000000d00cc3400000000000000000000000000000000000000000c00d00000000000000000000000000000000000000000000c00100100000000000000000000000000000000000000000c00400100000000000000000000000000000000000000000c00700100000000000000000000000000000000000000000c00a00100000000000000000000000000000000000000000c00d00100000000000000000000000000000000000000000c00000200000000000000000000000000000000000000000c00300200000000000000000000000000000000000000000c00800200000000000000000000000000000000000000000d00784b00000000000000000000000000000000000000000d00e53000000000000000000000000000000000000000000c00b00200000000000000000000000000000000000000000c00e00200000000000000000000000000000000000000000c00100300000000000000000000000000000000000000000c00400300000000000000000000000000000000000000000c00700300000000000000000000000000000000000000000c00a00300000000000000000000000000000000000000000c00d00300000000000000000000000000000000000000000c00000400000000000000000000000000000000000000000c00300400000000000000000000000000000000000000000c00800400000000000000000000000000000000000000000c00b00400000000000000000000000000000000000000000c00000500000000000000000000000000000000000000000c00300500000000000000000000000000000000000000000c00800500000000000000000000000000000000000000000c00b00500000000000000000000000000000000000000000c00f00500000000000000000000000000000000000000000c00600600000000000000000000000000000000000000000c00b00600000000000000000000000000000000000000000c00f00600000000000000000000000000000000000000000c00200700000000000000000000000000000000000000000c00500700000000000000000000000000000000000000000d008b3b00000000000000000000000000000000000000000d00043000000000000000000000000000000000000000000d00981800000000000000000000000000000000000000000d003d2d00000000000000000000000000000000000000000d00123400000000000000000000000000000000000000000d001d2b00000000000000000000000000000000000000000d00c12800000000000000000000000000000000000000000d00ea1d00000000000000000000000000000000000000000d00db0700000000000000000000000000000000000000000d00fe2400000000000000000000000000000000000000000d00c51b00000000000000000000000000000000000000000d00591800000000000000000000000000000000000000000d00e73100000000000000000000000000000000000000000d00ed3100000000000000000000000000000000000000000d00874d00000000000000000000000000000000000000000d007f1b00000000000000000000000000000000000000000d00ac0900000000000000000000000000000000000000000d00434d00000000000000000000000000000000000000000d00171000000000000000000000000000000000000000000d00d10900000000000000000000000000000000000000000d00943c00000000000000000000000000000000000000000c00800700000000000000000000000000000000000000000c00b00700000000000000000000000000000000000000000c00e00700000000000000000000000000000000000000000c00100800000000000000000000000000000000000000000c00400800000000000000000000000000000000000000000c00700800000000000000000000000000000000000000000c00a00800000000000000000000000000000000000000000c00e00800000000000000000000000000000000000000000d00f10100000000000000000000000000000000000000000d00244000000000000000000000000000000000000000000d000c3c00000000000000000000000000000000000000000d003b3b00000000000000000000000000000000000000000d007e3800000000000000000000000000000000000000000c00100a00000000000000000000000000000000000000000c00400a00000000000000000000000000000000000000000c00700a00000000000000000000000000000000000000000c00a00a00000000000000000000000000000000000000000c00d00a00000000000000000000000000000000000000000c00000b00000000000000000000000000000000000000000d00b14000000000000000000000000000000000000000000d00454800000000000000000000000000000000000000000d00920400000000000000000000000000000000000000000d003d1b00000000000000000000000000000000000000000d00a32400000000000000000000000000000000000000000d00432b00000000000000000000000000000000000000000d00474d00000000000000000000000000000000000000000d00664a00000000000000000000000000000000000000000d006f0a00000000000000000000000000000000000000000c00b00b00000000000000000000000000000000000000000c00e00b00000000000000000000000000000000000000000c00100c00000000000000000000000000000000000000000c00400c00000000000000000000000000000000000000000c00700c00000000000000000000000000000000000000000c00b00c00000000000000000000000000000000000000000d00641e00000000000000000000000000000000000000000d006d4b00000000000000000000000000000000000000000d00291e00000000000000000000000000000000000000000d000f3000000000000000000000000000000000000000000d00a30900000000000000000000000000000000000000000d000b3800000000000000000000000000000000000000000d00321b00000000000000000000000000000000000000000d00143000000000000000000000000000000000000000000d00ec0400000000000000000000000000000000000000000d00cf0e00000000000000000000000000000000000000000d00114d00000000000000000000000000000000000000000d00503000000000000000000000000000000000000000000d00dc3a00000000000000000000000000000000000000000d004b0500000000000000000000000000000000000000000c00f00c00000000000000000000000000000000000000000c00200d00000000000000000000000000000000000000000c00500d00000000000000000000000000000000000000000c00800d00000000000000000000000000000000000000000c00b00d00000000000000000000000000000000000000000c00e00d00000000000000000000000000000000000000000d00553400000000000000000000000000000000000000000d00932400000000000000000000000000000000000000000d00d43200000000000000000000000000000000000000000c00300b00000000000000000000000000000000000000000d00ae1900000000000000000000000000000000000000000d00da3200000000000000000000000000000000000000000d00144800000000000000000000000000000000000000000d00514f00000000000000000000000000000000000000000d00a74b00000000000000000000000000000000000000000d00774500000000000000000000000000000000000000000d00a24500000000000000000000000000000000000000000c00700b00000000000000000000000000000000000000000d00e53a00000000000000000000000000000000000000000d002a0a00000000000000000000000000000000000000000d00da1000000000000000000000000000000000000000000d00d30c00000000000000000000000000000000000000000d004b3300000000000000000000000000000000000000000d00251100000000000000000000000000000000000000000d00db3c00000000000000000000000000000000000000000d00ce4d00000000000000000000000000000000000000000d004d4c00000000000000000000000000000000000000000d00340a00000000000000000000000000000000000000000d00b54f00000000000000000000000000000000000000000d00242f00000000000000000000000000000000000000000d00d00700000000000000000000000000000000000000000d002a2f00000000000000000000000000000000000000000d00b01000000000000000000000000000000000000000000d00df3c00000000000000000000000000000000000000000d00ab0a00000000000000000000000000000000000000000d008e1100000000000000000000000000000000000000000d009d3400000000000000000000000000000000000000000d00a11e00000000000000000000000000000000000000000d00202500000000000000000000000000000000000000000d00663600000000000000000000000000000000000000000d000e4900000000000000000000000000000000000000000d00153e00000000000000000000000000000000000000000d00c10100000000000000000000000000000000000000000d00712c00000000000000000000000000000000000000000d00764400000000000000000000000000000000000000000d006b4e00000000000000000000000000000000000000000d005a4100000000000000000000000000000000000000000d00a01c00000000000000000000000000000000000000000d00064000000000000000000000000000000000000000000d00383900000000000000000000000000000000000000000d00120000000000000000000000000000000000000000000d00a41b00000000000000000000000000000000000000000d00812f00000000000000000000000000000000000000000d00094d00000000000000000000000000000000000000000d00e13400000000000000000000000000000000000000000d007c2300000000000000000000000000000000000000000d008c2300000000000000000000000000000000000000000d004b3700000000000000000000000000000000000000000d00614e00000000000000000000000000000000000000000d00ef3900000000000000000000000000000000000000000d00740b00000000000000000000000000000000000000000d00ff3d00000000000000000000000000000000000000000d004d0c00000000000000000000000000000000000000000d001a1d00000000000000000000000000000000000000000d002c4500000000000000000000000000000000000000000d008a1200000000000000000000000000000000000000000d00d11b00000000000000000000000000000000000000000d00501c00000000000000000000000000000000000000000d00fc2900000000000000000000000000000000000000000d00404700000000000000000000000000000000000000000d009a4a00000000000000000000000000000000000000000d002c2700000000000000000000000000000000000000000d00fb4000000000000000000000000000000000000000000d00180600000000000000000000000000000000000000000d00124100000000000000000000000000000000000000000d00924400000000000000000000000000000000000000000d00620900000000000000000000000000000000000000000d003a2a00000000000000000000000000000000000000000d00862a00000000000000000000000000000000000000000d00443b00000000000000000000000000000000000000000d00ee3d00000000000000000000000000000000000000000d00b41a00000000000000000000000000000000000000000d00d11200000000000000000000000000000000000000000d00e64400000000000000000000000000000000000000000d002f3200000000000000000000000000000000000000000d00c62700000000000000000000000000000000000000000d00da0900000000000000000000000000000000000000000d005b0e00000000000000000000000000000000000000000d002b1900000000000000000000000000000000000000000d004c0400000000000000000000000000000000000000000d000a1b00000000000000000000000000000000000000000d00b60700000000000000000000000000000000000000000d00fa4500000000000000000000000000000000000000000d00c93c00000000000000000000000000000000000000000d00b40300000000000000000000000000000000000000000d00af0500000000000000000000000000000000000000000d00d93400000000000000000000000000000000000000000d00613700000000000000000000000000000000000000000d00f62a00000000000000000000000000000000000000000d00f20d00000000000000000000000000000000000000000d00ff1200000000000000000000000000000000000000000d00844100000000000000000000000000000000000000000d00fe3300000000000000000000000000000000000000000d00793a00000000000000000000000000000000000000000d00fa0100000000000000000000000000000000000000000d00ee4900000000000000000000000000000000000000000d00403200000000000000000000000000000000000000000d00cd1800000000000000000000000000000000000000000d00e91500000000000000000000000000000000000000000d009e0d00000000000000000000000000000000000000000d00801500000000000000000000000000000000000000000d00e73e00000000000000000000000000000000000000000d005e1d00000000000000000000000000000000000000000d00a64000000000000000000000000000000000000000000d00083000000000000000000000000000000000000000000d00391900000000000000000000000000000000000000000d00f53e00000000000000000000000000000000000000000d002d3f00000000000000000000000000000000000000000d002c4b00000000000000000000000000000000000000000d00db1d00000000000000000000000000000000000000000d00721000000000000000000000000000000000000000000d00f84100000000000000000000000000000000000000000d007a2f00000000000000000000000000000000000000000d00b62b00000000000000000000000000000000000000000d00984600000000000000000000000000000000000000000d005e1300000000000000000000000000000000000000000d002b2500000000000000000000000000000000000000000d00b53f00000000000000000000000000000000000000000d00fc4200000000000000000000000000000000000000000d007b3900000000000000000000000000000000000000000d00f60000000000000000000000000000000000000000000d00ec0800000000000000000000000000000000000000000d00b60f00000000000000000000000000000000000000000d00a61100000000000000000000000000000000000000000d00ac1100000000000000000000000000000000000000000d00602900000000000000000000000000000000000000000d00ea3c00000000000000000000000000000000000000000d00670d00000000000000000000000000000000000000000d00cf4300000000000000000000000000000000000000000d00b61100000000000000000000000000000000000000000d00704a00000000000000000000000000000000000000000d005d3100000000000000000000000000000000000000000d00613100000000000000000000000000000000000000000d00a61e00000000000000000000000000000000000000000d00e84d00000000000000000000000000000000000000000d00ad4600000000000000000000000000000000000000000d00c32000000000000000000000000000000000000000000d00e14d00000000000000000000000000000000000000000d002b0800000000000000000000000000000000000000000d009e1300000000000000000000000000000000000000000d000c0000000000000000000000000000000000000000000d00174900000000000000000000000000000000000000000d00a51700000000000000000000000000000000000000000d00590000000000000000000000000000000000000000000d00961c00000000000000000000000000000000000000000d00630600000000000000000000000000000000000000000d00822700000000000000000000000000000000000000000d006c1400000000000000000000000000000000000000000d00d32300000000000000000000000000000000000000000d00df0800000000000000000000000000000000000000000d004b4900000000000000000000000000000000000000000d00712200000000000000000000000000000000000000000d00844a00000000000000000000000000000000000000000d00822200000000000000000000000000000000000000000d00080000000000000000000000000000000000000000000d00280b00000000000000000000000000000000000000000d008c1b00000000000000000000000000000000000000000d00230f00000000000000000000000000000000000000000d00a14600000000000000000000000000000000000000000d00652000000000000000000000000000000000000000000d002b0900000000000000000000000000000000000000000d00a51a00000000000000000000000000000000000000000d001f4100000000000000000000000000000000000000000d00231400000000000000000000000000000000000000000d002a2c00000000000000000000000000000000000000000d00d20100000000000000000000000000000000000000000d00584c00000000000000000000000000000000000000000d00f14d00000000000000000000000000000000000000000d001f0100000000000000000000000000000000000000000d00da1b00000000000000000000000000000000000000000d00bb3200000000000000000000000000000000000000000d00172800000000000000000000000000000000000000000d00620c00000000000000000000000000000000000000000d005a4500000000000000000000000000000000000000000d00e82d00000000000000000000000000000000000000000d00c93200000000000000000000000000000000000000000d00680b00000000000000000000000000000000000000000d00ba4000000000000000000000000000000000000000000d00f43f00000000000000000000000000000000000000000d00bf2b00000000000000000000000000000000000000000d00c23900000000000000000000000000000000000000000d00d80f00000000000000000000000000000000000000000d00fe2b00000000000000000000000000000000000000000d00172300000000000000000000000000000000000000000d00592300000000000000000000000000000000000000000d003d3900000000000000000000000000000000000000000d00e33600000000000000000000000000000000000000000d00b62900000000000000000000000000000000000000000d008d4a00000000000000000000000000000000000000000d00a80d00000000000000000000000000000000000000000d000e2c00000000000000000000000000000000000000000d00e93600000000000000000000000000000000000000000d00253700000000000000000000000000000000000000000d000a0400000000000000000000000000000000000000000d00964000000000000000000000000000000000000000000d00a73300000000000000000000000000000000000000000d00240100000000000000000000000000000000000000000d00ab0500000000000000000000000000000000000000000d00174b00000000000000000000000000000000000000000d00e54e00000000000000000000000000000000000000000d001f4b00000000000000000000000000000000000000000d00652800000000000000000000000000000000000000000d006a2e00000000000000000000000000000000000000000d00263500000000000000000000000000000000000000000d00204900000000000000000000000000000000000000000d00b63d00000000000000000000000000000000000000000d00b71b00000000000000000000000000000000000000000d00a33400000000000000000000000000000000000000000d00570f00000000000000000000000000000000000000000d00822d00000000000000000000000000000000000000000d006a1500000000000000000000000000000000000000000d00bd4700000000000000000000000000000000000000000d00bb4a00000000000000000000000000000000000000000d00a20d00000000000000000000000000000000000000000d00ec0000000000000000000000000000000000000000000d00401a00000000000000000000000000000000000000000d00e03600000000000000000000000000000000000000000d008a2400000000000000000000000000000000000000000d00233c00000000000000000000000000000000000000000d00342b00000000000000000000000000000000000000000d00954700000000000000000000000000000000000000000d00f63100000000000000000000000000000000000000000d006b3a00000000000000000000000000000000000000000d001a4d00000000000000000000000000000000000000000d001f2c00000000000000000000000000000000000000000d007e0900000000000000000000000000000000000000000d00e50800000000000000000000000000000000000000000d00a03300000000000000000000000000000000000000000d00790f00000000000000000000000000000000000000000d009c0500000000000000000000000000000000000000000d00034700000000000000000000000000000000000000000d00df3d00000000000000000000000000000000000000000d00ba0300000000000000000000000000000000000000000d00824400000000000000000000000000000000000000000d00f60600000000000000000000000000000000000000000d00a70e00000000000000000000000000000000000000000d007b4200000000000000000000000000000000000000000d00bb3c00000000000000000000000000000000000000000d00bc2f00000000000000000000000000000000000000000d00ae4a00000000000000000000000000000000000000000d001e4a00000000000000000000000000000000000000000d00444f00000000000000000000000000000000000000000d00ec2a00000000000000000000000000000000000000000d002d1700000000000000000000000000000000000000000d00e93000000000000000000000000000000000000000000d00604000000000000000000000000000000000000000000d00091300000000000000000000000000000000000000000d00411000000000000000000000000000000000000000000d004b3400000000000000000000000000000000000000000d00103300000000000000000000000000000000000000000d00644500000000000000000000000000000000000000000d00051b00000000000000000000000000000000000000000d00bc2700000000000000000000000000000000000000000d00554800000000000000000000000000000000000000000d001c3500000000000000000000000000000000000000000d00c20200000000000000000000000000000000000000000d00fa1400000000000000000000000000000000000000000d00180500000000000000000000000000000000000000000d001d1300000000000000000000000000000000000000000d00664b00000000000000000000000000000000000000000d00313500000000000000000000000000000000000000000d00e11900000000000000000000000000000000000000000d00320700000000000000000000000000000000000000000d00823a00000000000000000000000000000000000000000d00740700000000000000000000000000000000000000000d003a3f00000000000000000000000000000000000000000d00063300000000000000000000000000000000000000000d000b4200000000000000000000000000000000000000000d000d0a00000000000000000000000000000000000000000d00112800000000000000000000000000000000000000000d00211900000000000000000000000000000000000000000d000a2400000000000000000000000000000000000000000d008f2d00000000000000000000000000000000000000000d002d1100000000000000000000000000000000000000000c00f00f00000000000000000000000000000000000000000c00201000000000000000000000000000000000000000000c00501000000000000000000000000000000000000000000d00f10600000000000000000000000000000000000000000d00033800000000000000000000000000000000000000000d00e12e00000000000000000000000000000000000000000d006a1900000000000000000000000000000000000000000d00731900000000000000000000000000000000000000000d00142f00000000000000000000000000000000000000000d00721600000000000000000000000000000000000000000d00084800000000000000000000000000000000000000000400406e010000000000000000000000000000000000000004004e6e010000000000000000000000000000000000000004002eb30100000000000000000000000000000000000000040030b30100000000000000000000000000000000000000040072b40100000000000000000000000000000000000000040056b601000000000000000000000000000000000000000400acb60100000000000000000000000000000000000000040024ba0100000000000000000000000000000000000000040032ba01000000000000000000000000000000000000000400b0bb01000000000000000000000000000000000000000400c2bb01000000000000000000000000000000000000000400d4bb01000000000000000000000000000000000000000400e2bb01000000000000000000000000000000000000000400f0bb01000000000000000000000000000000000000000400febb010000000000000000000000000000000000000004006ebc010000000000000000000000000000000000000004002abe01000000000000000000000000000000000000000400debe0100000000000000000000000000000000000000040016bf0100000000000000000000000000000000000000040020bf01000000000000000000000000000000000000000400d6bf0100000000000000000000000000000000000000040010c00100000000000000000000000000000000000000040030c10100000000000000000000000000000000000000040030c201000000000000000000000000000000000000000400c8c201000000000000000000000000000000000000000400d6c20100000000000000000000000000000000000000040048c301000000000000000000000000000000000000000400bac301000000000000000000000000000000000000000400d0c30100000000000000000000000000000000000000040072c401000000000000000000000000000000000000000400e2c401000000000000000000000000005a6900000400f1ff00000000000000000000000000000000686900000200040092940200000000003e000000000000006f69000000000400929402000000000000000000000000007269000002000400d0940200000000000e000000000000008569000000000400d0940200000000000000000000000000886900000100070098ca02000000000008000000000000009369000002000400de94020000000000c21a000000000000a469000000000400de940200000000000000000000000000a769000002000400a0af020000000000ae00000000000000bd69000000000400a0af0200000000000000000000000000c0690000000004004eb00200000000000000000000000000c369000000000400f0b00200000000000000000000000000c66900000000040042b10200000000000000000000000000c96900000000040058b10200000000000000000000000000cc69000000000400d2940200000000000000000000000000d1690000000004002c950200000000000000000000000000d66900000000040040950200000000000000000000000000db6900000000040088950200000000000000000000000000e0690000000004009a950200000000000000000000000000e569000000000400ec950200000000000000000000000000ea69000000000400f4950200000000000000000000000000ef6900000000040046960200000000000000000000000000f46900000000040050960200000000000000000000000000f96900000000040004950200000000000000000000000000fd690000000004006caf0200000000000000000000000000016a0000000004000cb00200000000000000000000000000066a00000000040030b002000000000000000000000000000b6a00000000040002b00200000000000000000000000000106a0000000004006cb00200000000000000000000000000156a00000000040076b002000000000000000000000000001a6a00000000040080b002000000000000000000000000001f6a0000000004008ab00200000000000000000000000000246a00000000040094b00200000000000000000000000000296a0000000004009eb002000000000000000000000000002e6a000000000400a8b00200000000000000000000000000336a000000000400b2b00200000000000000000000000000386a000000000400c2b002000000000000000000000000003d6a00000000040034b10200000000000000000000000000426a00000000040054b10200000000000000000000000000476a00000000040024b202000000000000000000000000004c6a000000000400a2b10200000000000000000000000000516a000000000400cab10200000000000000000000000000566a00000400f1ff000000000000000000000000000000005c6a00000000040030b202000000000000000000000000005f6a000000000400feb20200000000000000000000000000626a00000000040026b70200000000000000000000000000656a0000000004004cb70200000000000000000000000000686a000000000400fcb202000000000000000000000000006c6a000000000400ecb20200000000000000000000000000706a00000000040022b70200000000000000000000000000756a000000000400dab302000000000000000000000000007a6a00000000040022b302000000000000000000000000007f6a000000000400c4b50200000000000000000000000000846a0000000004001eb30200000000000000000000000000896a000000000400eeb302000000000000000000000000008e6a0000000004009ab30200000000000000000000000000936a00000000040058b30200000000000000000000000000986a0000000004005cb602000000000000000000000000009d6a00000000040068b30200000000000000000000000000a26a000000000400c0b30200000000000000000000000000a76a000000000400ccb30200000000000000000000000000ac6a000000000400aeb50200000000000000000000000000b16a000000000400a2b40200000000000000000000000000b66a0000000004008cb60200000000000000000000000000bb6a000000000400ceb50200000000000000000000000000c06a00000000040038b40200000000000000000000000000c56a0000000004003cb50200000000000000000000000000ca6a00000000040084b50200000000000000000000000000cf6a000000000400aab50200000000000000000000000000d46a000000000400d0b30200000000000000000000000000d96a000000000400f0b50200000000000000000000000000de6a00000000040066b60200000000000000000000000000e36a000000000400b6b60200000000000000000000000000e86a00000000040036b30200000000000000000000000000ed6a0000000004003cb70200000000000000000000000000f36a00000000040040b70200000000000000000000000000f96a00000000040028b70200000000000000000000000000ff6a0000000004002cb80200000000000000000000000000056b0000000004000cb902000000000000000000000000000b6b00000000040030b80200000000000000000000000000116b00000000040098b80200000000000000000000000000176b00000000040012b902000000000000000000000000001d6b0000000004000eb90200000000000000000000000000236b000000000400aeb70200000000000000000000000000296b00000000040082b802000000000000000000000000002f6b00000000040028b90200000000000000000000000000356b0000000004004eb802000000000000000000000000003b6b00000000040048b80200000000000000000000000000416b00000000040018b90200000000000000000000000000476b0000000004006cb802000000000000000000000000004d6b0000000004002cb90200000000000000000000000000536b000000000400b0b80200000000000000000000000000596b000000000400aab802000000000000000000000000005f6b0000000004001cb90200000000000000000000000000656b000000000400d8b802000000000000000000000000006b6b000000000400fab80200000000000000000000000000716b000000000400f8b80200000000000000000000000000776b000000000400f4b802000000000000000000000000007d6b00000000040062b80200000000000000000000000000836b000000000400c2b802000000000000000000000000009f6b0000020204004cb7020000000000e601000000000000a76b000002020400feb20200000000002804000000000000ae6b00000202040026b70200000000002600000000000000b56b00000202040030b2020000000000ce00000000000000896b000012000400e0470100000000009025000000000000986b00001000040074360100000000000000000000000000bc6b00001200040042b10200000000001600000000000000cb6b00001200040058b1020000000000d800000000000000d96b000012000400f0b00200000000005200000000000000f56b0000120004004eb0020000000000a200000000000000002e726f64617461002e73726f646174612e63737438002e65685f6672616d65002e74657874002e7364617461002e64617461002e73646174612e6d656d7365745f762e30002e627373002e64656275675f616262726576002e64656275675f696e666f002e64656275675f6172616e676573002e64656275675f72616e676573002e64656275675f737472002e64656275675f7075626e616d6573002e64656275675f7075627479706573002e72697363762e61747472696275746573002e64656275675f6c696e65002e636f6d6d656e74002e73796d746162002e7368737472746162002e73747274616200007374616b655f736d742e646436616664343835633633343335632d6367752e30002e4c435049305f30005f5a4e34636f72653370747231373364726f705f696e5f706c616365244c5424616c6c6f632e2e7665632e2e696e746f5f697465722e2e496e746f49746572244c5424244c502424753562247538247533622424753230243230247535642424432424753562247538247533622424753230243332247535642424432461786f6e5f74797065732e2e67656e6572617465642e2e7374616b655f7265616465722e2e5374616b65496e666f44656c74612452502424475424244754243137683236336137653365303866636139333745002e4c706372656c5f686930005f5a4e36345f244c5424616c6c6f632e2e72632e2e5263244c54245424475424247532302461732475323024636f72652e2e6f70732e2e64726f702e2e44726f70244754243464726f703137683663346239333364656266363135663545005f5f727573745f6465616c6c6f63005f5a4e34636f726533707472343664726f705f696e5f706c616365244c5424616c6c6f632e2e7665632e2e566563244c5424753824475424244754243137683361313733353239636533623265663445005f5a4e34636f726533707472383864726f705f696e5f706c616365244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e7365742e2e4254726565536574244c54247574696c2e2e736d742e2e4c6f636b496e666f24475424244754243137683665343465643866393463343166666345002e4c706372656c5f686931002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e30005f5a4e34636f72653970616e69636b696e673570616e69633137686437373538656430613265383739363145005f5a4e35616c6c6f633131636f6c6c656374696f6e733562747265653373657432314254726565536574244c542454244324412447542436696e736572743137686464393035633939376636373034323545005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565367365617263683134325f244c5424696d706c2475323024616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e4e6f6465526566244c5424426f72726f77547970652443244b24432456244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4c6561664f72496e7465726e616c244754242447542431317365617263685f747265653137683334313732383863663534343435313045005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f646532314c6561664e6f6465244c54244b2443245624475424336e65773137683030343135616633666232326365633045005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f64653235496e7465726e616c4e6f6465244c54244b2443245624475424336e65773137683032323863313432336565363266306545005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f646532313448616e646c65244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e4e6f6465526566244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4d75742443244b24432456244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e496e7465726e616c24475424244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e45646765244754243130696e736572745f6669743137686333643836376265346235366332393945002e4c706372656c5f686934002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3639002e4c706372656c5f686935002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3635005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243135636f70795f66726f6d5f736c69636531376c656e5f6d69736d617463685f6661696c3137686531663934356265353831313135613845002e4c706372656c5f686936002e4c706372656c5f686932002e4c706372656c5f686933002e4c706372656c5f686937002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3537002e4c706372656c5f686938005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f64653132354e6f6465526566244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4d75742443244b24432456244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4c6561664f72496e7465726e616c24475424313663686f6f73655f706172656e745f6b763137683139343665383636343762653264393545005f5a4e34636f72653970616e69636b696e67313870616e69635f6e6f756e77696e645f666d743137683133386130386530383963323036303445005f5f727573745f616c6c6f63005f5f727573745f616c6c6f635f6572726f725f68616e646c6572005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b2443245624475424313562756c6b5f737465616c5f6c6566743137686539616634316334303135636434623645002e4c706372656c5f686939002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3733002e4c706372656c5f68693131002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3735002e4c706372656c5f68693130002e4c706372656c5f68693132002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3737005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b2443245624475424313662756c6b5f737465616c5f72696768743137686162393832373662656263346330393645002e4c706372656c5f68693133002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3830002e4c706372656c5f68693135002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3832002e4c706372656c5f68693134002e4c706372656c5f68693136005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b244324562447542432356d657267655f747261636b696e675f6368696c645f656467653137683538306266633666353961646136383045002e4c706372656c5f68693138002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3835002e4c706372656c5f68693137002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3837005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b244324562447542438646f5f6d657267653137683762346633316135393139303638643245002e4c706372656c5f68693139005f5a4e35616c6c6f633131636f6c6c656374696f6e733562747265653672656d6f76653235395f244c5424696d706c2475323024616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e48616e646c65244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e4e6f6465526566244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4d75742443244b24432456244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4c65616624475424244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4b562447542424475424313472656d6f76655f6c6561665f6b763137683034323333323932386162316238636645002e4c706372656c5f68693230005f5a4e37636b625f73746433656e7634415247563137683036373561626564353032343439613545005f5a4e37636b625f7374643130686967685f6c6576656c31316c6f61645f7363726970743137683962326234613433643962613162666545005f5a4e3131636b625f747970655f696431366861735f747970655f69645f63656c6c3137683163316466616433653431643434383645005f5a4e38345f244c54247574696c2e2e6572726f722e2e4572726f72247532302461732475323024636f72652e2e636f6e766572742e2e46726f6d244c5424636b625f747970655f69642e2e4572726f7224475424244754243466726f6d3137683537363538306531656461613935643645005f5a4e347574696c3668656c706572313663616c635f7363726970745f686173683137686361393462346333346566393134393545005f5a4e35616c6c6f63377261775f7665633139526177566563244c54245424432441244754243131616c6c6f636174655f696e3137683961373435623837316432623838663945005f5a4e347574696c3668656c70657232376765745f63656c6c5f636f756e745f62795f747970655f686173683137683636366663636666636434353161366445005f5a4e37636b625f7374643130686967685f6c6576656c31396c6f61645f63656c6c5f747970655f686173683137686661353738353337303831333261613945005f5a4e39305f244c54247574696c2e2e6572726f722e2e4572726f72247532302461732475323024636f72652e2e636f6e766572742e2e46726f6d244c5424636b625f7374642e2e6572726f722e2e5379734572726f7224475424244754243466726f6d3137686233643163343538633564356263343545002e4c706372656c5f68693234002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e383436002e4c706372656c5f68693236005f5a4e37636b625f7374643130686967685f6c6576656c31306c6f61645f696e7075743137686333316231653162623031363962653245002e4c706372656c5f68693233005f5a4e3130626c616b6532625f727337626c616b6532623134426c616b6532624275696c646572356275696c643137683463643438663738663037316532306145002e4c706372656c5f68693235005f5a4e34636f726533707472353564726f705f696e5f706c616365244c54246d6f6c6563756c652e2e6572726f722e2e566572696669636174696f6e4572726f72244754243137683936383830623737653965663033383845002e4c706372656c5f68693237002e4c706372656c5f68693238002e4c706372656c5f68693239002e4c706372656c5f68693231007374722e342e3733005f5a4e34636f726535736c69636535696e64657837345f244c5424696d706c2475323024636f72652e2e6f70732e2e696e6465782e2e496e646578244c542449244754242475323024666f72247532302424753562245424753564242447542435696e6465783137683064326565363561653136626361336545005f5a4e3131315f244c5424616c6c6f632e2e7665632e2e566563244c54245424475424247532302461732475323024616c6c6f632e2e7665632e2e737065635f66726f6d5f697465725f6e65737465642e2e5370656346726f6d497465724e6573746564244c5424542443244924475424244754243966726f6d5f697465723137683032353562336632346332623633633445005f5a4e35616c6c6f63337665633136566563244c542454244324412447542434707573683137683832346530366138613965323339383745005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f7233616e793137683031323866356465313834336464653445002e4c706372656c5f68693331002e4c706372656c5f68693232007374722e302e313130002e4c706372656c5f68693330005f5a4e3130325f244c5424636b625f7374616e64616c6f6e655f74797065732e2e67656e6572617465642e2e626c6f636b636861696e2e2e42797465735265616465722475323024617324753230246d6f6c6563756c652e2e7072656c7564652e2e52656164657224475424367665726966793137683135663233383466353032373265326345005f5a4e386d6f6c6563756c6535627974657335427974657335736c6963653137683133633337653065643765643238336345005f5a4e3230636b625f7374616e64616c6f6e655f74797065733967656e6572617465643130626c6f636b636861696e354279746573387261775f646174613137686165613062386538653731396665363945005f5a4e347574696c3668656c70657231386765745f7374616b655f736d745f646174613137683531393538393938623361383432363145005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231365374616b65536d7443656c6c4461746131366d657461646174615f747970655f69643137683333316537333761333766666465306145005f5a4e347574696c3668656c70657231326765745f747970655f6964733137683161323938396534376363663639393545005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f72656164657237547970654964733134787564745f747970655f686173683137686334653636633566343738343237356145005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f726561646572375479706549647331397374616b655f736d745f636f64655f686173683137683939313230643232643561376161363745005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f726561646572375479706549647331377374616b655f736d745f747970655f69643137683133613730383736373561386135323245005f5a4e347574696c3668656c70657231356765745f7363726970745f686173683137683861333134336361336163636135633445005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f72656164657237547970654964733230636865636b706f696e745f636f64655f686173683137683561366363373337366465333564383045005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f72656164657237547970654964733138636865636b706f696e745f747970655f69643137683062376537323033303666383865346345005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f7265616465723754797065496473313877697468647261775f636f64655f686173683137686636356461336666633664366137323445005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f726561646572375479706549647331386d657461646174615f636f64655f686173683137683263623137613437626166656264306645005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f726561646572375479706549647331366d657461646174615f747970655f69643137683833306539326563613930383864363745005f5a4e3230636b625f7374616e64616c6f6e655f74797065733967656e6572617465643130626c6f636b636861696e31315769746e65737341726773346c6f636b3137686233326333343036613431316531636245005f5a4e39385f244c54246d6f6c6563756c65322e2e7265616465722e2e437572736f72247532302461732475323024636f72652e2e636f6e766572742e2e46726f6d244c5424616c6c6f632e2e7665632e2e566563244c542475382447542424475424244754243466726f6d3137686365383937663564613837343036643045005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231345374616b65496e666f44656c7461313169735f696e6372656173653137683166386136356661303836623163316645005f5a4e347574696c3668656c70657231376765745f63757272656e745f65706f63683137683433313039626562306665666534313945005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231385374616b65536d74557064617465496e666f3135616c6c5f7374616b655f696e666f733137686331656532343334363962343463366245005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231305374616b65496e666f73336c656e3137683862303137666338646362303233393945005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231305374616b65496e666f73336765743137683536663765343736643831623335613045005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f726561646572395374616b65496e666f34616464723137683737663935343236353164653934373045005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231345374616b65496e666f44656c746136616d6f756e743137683736303137613463316430633135626445005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231385374616b65536d74557064617465496e666f31356f6c645f65706f63685f70726f6f663137683835396638343561623737663561346545005f5a4e347574696c33736d7431317536345f746f5f683235363137683630616266646338653134653935363145005f5a4e347574696c33736d7431377665726966795f326c617965725f736d743137683133343062636139316137313632616545005f5a4e347574696c3668656c70657232326765745f7374616b655f7570646174655f696e666f733137686337343437303336323761616365383045005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231345374616b65496e666f44656c74613138696e61756775726174696f6e5f65706f63683137683538323561303933383837366165313345005f5a4e347574696c3668656c70657233306765745f7374616b655f61745f646174615f62795f6c6f636b5f686173683137683536356232313136353933333665623945005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231355374616b65417443656c6c446174613564656c74613137683762333332613765343438316530613845005f5a4e3130385f244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6d61702e2e49746572244c54244b2443245624475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683932393561376437613164316266393145005f5a4e347574696c3668656c706572323563616c635f7769746864726177616c5f6c6f636b5f686173683137683038613966633761623133353165326345005f5a4e347574696c3668656c70657233336765745f77697468647261775f61745f646174615f62795f6c6f636b5f686173683137686531356438613763623138663661663445005f5a4e347574696c3668656c70657231356765745f71756f72756d5f73697a653137683930353932376137656234333038306645005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231385374616b65536d74557064617465496e666f31356e65775f65706f63685f70726f6f663137686236623761343265306435646564653745002e4c706372656c5f68693332002e4c706372656c5f68693433007374722e31002e4c706372656c5f68693333002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3436002e4c706372656c5f68693334002e4c616e6f6e2e36633237623166666234666234346562313164656530663863336331326232322e33005f5a4e34636f726536726573756c743133756e777261705f6661696c65643137683030653934303161326339653536633045002e4c706372656c5f68693435002e4c706372656c5f68693436002e4c706372656c5f68693335002e4c706372656c5f68693336002e4c616e6f6e2e36633237623166666234666234346562313164656530663863336331326232322e32002e4c706372656c5f68693337002e4c706372656c5f68693338002e4c706372656c5f68693339002e4c706372656c5f68693430002e4c706372656c5f68693431002e4c706372656c5f68693432002e4c706372656c5f68693434002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e363300727573745f626567696e5f756e77696e64005f5a4e37636b625f7374643873797363616c6c73366e617469766534657869743137683163616638653234666532613530323145005f5f72675f616c6c6f63005f5a4e3130365f244c542462756464795f616c6c6f632e2e6e6f6e5f746872656164736166655f616c6c6f632e2e4e6f6e54687265616473616665416c6c6f63247532302461732475323024636f72652e2e616c6c6f632e2e676c6f62616c2e2e476c6f62616c416c6c6f632447542435616c6c6f633137683966656332343337626566343266383945005f5f72675f6465616c6c6f63005f5a4e3130365f244c542462756464795f616c6c6f632e2e6e6f6e5f746872656164736166655f616c6c6f632e2e4e6f6e54687265616473616665416c6c6f63247532302461732475323024636f72652e2e616c6c6f632e2e676c6f62616c2e2e476c6f62616c416c6c6f6324475424376465616c6c6f633137686530336235656339643238613732396445005f5f72675f7265616c6c6f63005f5f72675f616c6c6f635f7a65726f6564005f5f727573745f7265616c6c6f63005f5f727573745f616c6c6f635f7a65726f6564005f5f72646c5f6f6f6d005f5a4e35616c6c6f63377261775f766563313763617061636974795f6f766572666c6f773137683736396433373734353939336431626545005f5a4e396d6f6c6563756c65323672656164657236437572736f72323164796e7665635f736c6963655f62795f696e6465783137683464633230383535323662653634303045005f5a4e396d6f6c6563756c6532367265616465723130385f244c5424696d706c2475323024636f72652e2e636f6e766572742e2e46726f6d244c54246d6f6c6563756c65322e2e7265616465722e2e437572736f72244754242475323024666f722475323024616c6c6f632e2e7665632e2e566563244c5424753824475424244754243466726f6d3137683965653331373661666261663535343545002e4c706372656c5f68693437002e4c706372656c5f68693438002e4c616e6f6e2e65383134633736363361666663333138633766356639363865643531663662352e3139002e4c706372656c5f68693439002e4c706372656c5f68693530002e4c706372656c5f68693531002e4c706372656c5f68693532002e4c706372656c5f68693533002e4c706372656c5f68693534002e4c706372656c5f68693535002e4c706372656c5f68693536002e4c706372656c5f68693537002e4c706372656c5f68693538002e4c706372656c5f68693539002e4c706372656c5f68693630002e4c706372656c5f68693631002e4c706372656c5f68693632005f5a4e396d6f6c6563756c65323672656164657238355f244c5424696d706c2475323024636f72652e2e636f6e766572742e2e46726f6d244c54246d6f6c6563756c65322e2e7265616465722e2e437572736f72244754242475323024666f7224753230247538244754243466726f6d3137686461653235633931336631613435396545002e4c706372656c5f68693633002e4c706372656c5f68693634002e4c706372656c5f68693635002e4c706372656c5f68693636005f5a4e396d6f6c6563756c65323672656164657238365f244c5424696d706c2475323024636f72652e2e636f6e766572742e2e46726f6d244c54246d6f6c6563756c65322e2e7265616465722e2e437572736f72244754242475323024666f722475323024753634244754243466726f6d3137686232663035653938653831303635333145002e4c706372656c5f68693637002e4c706372656c5f68693638002e4c706372656c5f68693639002e4c706372656c5f68693730002e4c706372656c5f68693731002e4c706372656c5f68693732002e4c706372656c5f68693733002e4c706372656c5f68693734005f5a4e396d6f6c6563756c65323672656164657236437572736f723876616c69646174653137683930306131623931383065653939313845005f5a4e396d6f6c6563756c65323672656164657236437572736f7231346765745f6974656d5f636f756e743137683362393033346337303939633162346445002e4c706372656c5f68693735002e4c706372656c5f68693736002e4c706372656c5f68693737002e4c706372656c5f68693738002e4c706372656c5f68693739002e4c706372656c5f68693830005f5a4e396d6f6c6563756c65323672656164657236437572736f723139636f6e766572745f746f5f72617762797465733137683634326263616436376665326537643145002e4c706372656c5f68693831002e4c706372656c5f68693832002e4c706372656c5f68693833002e4c706372656c5f68693834002e4c706372656c5f68693835002e4c706372656c5f68693836002e4c706372656c5f68693837002e4c706372656c5f68693838005f5a4e3131626c616b6532625f72656637777261707065723134426c616b6532624275696c646572356275696c643137683964636431366662373535323133626345005f5a4e3131626c616b6532625f7265663131626c616b6532625f7265663138626c616b6532625f696e69745f706172616d3137683431613831343963666239633164343445005f5a4e3131626c616b6532625f7265663131626c616b6532625f7265663134626c616b6532625f7570646174653137683337646637643338333264666265336545002e4c706372656c5f68693839005f5a4e3131626c616b6532625f7265663131626c616b6532625f7265663130626c616b6532625f49563137686532356438333932346363316638393145005f5a4e3131626c616b6532625f7265663131626c616b6532625f7265663136626c616b6532625f636f6d70726573733137683531363361326435303733336262323945002e4c43504934395f30002e4c43504934395f31002e4c43504934395f32002e4c43504934395f33002e4c43504934395f34002e4c43504934395f35002e4c43504934395f36002e4c43504934395f37002e4c706372656c5f68693930002e4c706372656c5f68693931002e4c706372656c5f68693932002e4c706372656c5f68693933002e4c706372656c5f68693934002e4c706372656c5f68693935002e4c706372656c5f68693936002e4c706372656c5f68693937005f5a4e3131626c616b6532625f726566377772617070657237426c616b6532623866696e616c697a653137683431356365303263316365386263623745005f5a4e313162756464795f616c6c6f63313162756464795f616c6c6f6331304275646479416c6c6f63336e65773137683039343964346234353436656265666245005f5a4e313162756464795f616c6c6f63313162756464795f616c6c6f6337726f756e6475703137686533656266373734346663663366363345002e4c706372656c5f6869313035007374722e342e3633005f5a4e313162756464795f616c6c6f63313162756464795f616c6c6f63366e626c6f636b3137683537623963376462363561386133343745005f5a4e313162756464795f616c6c6f63313162756464795f616c6c6f6331304275646479416c6c6f633131626c6f636b5f696e6465783137683333633165376336333564613363643945005f5a4e34636f7265366f7074696f6e31336578706563745f6661696c65643137686332333330616533386638616564396545002e4c706372656c5f6869313130002e4c706372656c5f6869313036002e4c706372656c5f6869313037002e4c706372656c5f68693938002e4c706372656c5f6869313030007374722e322e3634002e4c706372656c5f6869313031007374722e332e3635002e4c706372656c5f6869313032002e4c706372656c5f6869313033007374722e312e3632002e4c706372656c5f6869313034002e4c706372656c5f6869313131002e4c706372656c5f6869313038007374722e302e3631002e4c706372656c5f68693939002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3135002e4c706372656c5f6869313132002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3238005f5a4e34636f72653970616e69636b696e67313370616e69635f646973706c61793137683538303536323433613031393534316645002e4c706372656c5f6869313039002e4c706372656c5f6869313133002e4c706372656c5f6869313134002e4c706372656c5f6869313135002e4c706372656c5f6869313136002e4c706372656c5f6869313137002e4c706372656c5f6869313139002e4c706372656c5f6869313230002e4c706372656c5f6869313138002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3338005f5a4e313162756464795f616c6c6f633130666173745f616c6c6f633946617374416c6c6f63336e65773137683239303962396561363461333531383845002e4c706372656c5f6869313232002e4c706372656c5f6869313231002e4c706372656c5f6869313233002e4c706372656c5f6869313234005f5a4e397374616b655f736d7435414c4c4f433137683263336231343434623861633161633845002e4c706372656c5f6869313238002e4c706372656c5f6869313333002e4c706372656c5f6869313334002e4c706372656c5f6869313331002e4c706372656c5f6869313335002e4c706372656c5f6869313336002e4c706372656c5f6869313332002e4c706372656c5f6869313237002e4c706372656c5f6869313239002e4c706372656c5f6869313330002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e32002e4c706372656c5f6869313235002e4c706372656c5f6869313236002e4c706372656c5f6869313337002e4c706372656c5f6869313338002e4c706372656c5f6869313339002e4c706372656c5f6869313433002e4c706372656c5f6869313432002e4c706372656c5f6869313436002e4c706372656c5f6869313438002e4c706372656c5f6869313439002e4c706372656c5f6869313530002e4c706372656c5f6869313437002e4c706372656c5f6869313430002e4c706372656c5f6869313431002e4c706372656c5f6869313434002e4c706372656c5f6869313435005f5a4e35616c6c6f63377261775f7665633139526177566563244c54245424432441244754243131616c6c6f636174655f696e3137683334393639363464643031633234363645005f5a4e35616c6c6f63377261775f7665633139526177566563244c542454244324412447542437726573657276653231646f5f726573657276655f616e645f68616e646c653137686234636364626536643135363830353445002e4c706372656c5f6869313531007374722e302e3731005f5a4e35616c6c6f63377261775f7665633139526177566563244c5424542443244124475424313467726f775f616d6f7274697a65643137683131313435313531653037646531613245005f5a4e35616c6c6f63377261775f766563313166696e6973685f67726f773137683362363537323731663362336132663345005f5a4e35616c6c6f63377261775f7665633139526177566563244c54245424432441244754243136726573657276655f666f725f707573683137683364383734353931323332303230376445002e4c706372656c5f6869313532002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e313734002e4c706372656c5f6869313533002e4c706372656c5f6869313534005f5a4e3230636b625f7374616e64616c6f6e655f74797065733130636f6e76657273696f6e3130626c6f636b636861696e3134395f244c5424696d706c2475323024636b625f7374616e64616c6f6e655f74797065732e2e7072656c7564652e2e5061636b244c5424636b625f7374616e64616c6f6e655f74797065732e2e67656e6572617465642e2e626c6f636b636861696e2e2e427974653332244754242475323024666f72247532302424753562247538247533622424753230243332247535642424475424347061636b3137683838633365666265633136666335636345005f5a4e3230636b625f7374616e64616c6f6e655f74797065733130636f6e76657273696f6e397072696d69746976653133365f244c5424696d706c2475323024636b625f7374616e64616c6f6e655f74797065732e2e7072656c7564652e2e5061636b244c5424636b625f7374616e64616c6f6e655f74797065732e2e67656e6572617465642e2e626c6f636b636861696e2e2e4279746573244754242475323024666f72247532302424753562247538247535642424475424347061636b3137686534363231633861323935306563356145005f5a4e3133325f244c5424616c6c6f632e2e7665632e2e566563244c5424542443244124475424247532302461732475323024616c6c6f632e2e7665632e2e737065635f657874656e642e2e53706563457874656e64244c54242452462454244324636f72652e2e736c6963652e2e697465722e2e49746572244c5424542447542424475424244754243131737065635f657874656e643137683464663561353366366631653763336445002e4c706372656c5f6869313535007374722e322e3730005f5a4e39375f244c5424636b625f7374616e64616c6f6e655f74797065732e2e67656e6572617465642e2e626c6f636b636861696e2e2e5363726970742475323024617324753230246d6f6c6563756c652e2e7072656c7564652e2e456e746974792447542431316e65775f6275696c6465723137683663323863633439326130386634363645005f5a4e3130355f244c5424636b625f7374616e64616c6f6e655f74797065732e2e67656e6572617465642e2e626c6f636b636861696e2e2e5363726970744275696c6465722475323024617324753230246d6f6c6563756c652e2e7072656c7564652e2e4275696c64657224475424356275696c643137683462313334356436646334623638326145002e4c706372656c5f6869313536002e4c706372656c5f6869313537002e4c706372656c5f6869313538005f5a4e36315f244c5424636b625f7374642e2e6572726f722e2e5379734572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683863383033303266623836336136303845002e4c706372656c5f6869313539002e4c4a544937365f30002e4c424237365f31002e4c706372656c5f6869313630002e4c616e6f6e2e34313466363731613135666237623063306532636261396133343630323939342e3339002e4c424237365f32002e4c706372656c5f6869313631002e4c616e6f6e2e34313466363731613135666237623063306532636261396133343630323939342e3338002e4c424237365f33002e4c706372656c5f6869313632002e4c616e6f6e2e34313466363731613135666237623063306532636261396133343630323939342e3336002e4c706372656c5f6869313633002e4c616e6f6e2e34313466363731613135666237623063306532636261396133343630323939342e3337002e4c424237365f34002e4c706372656c5f6869313634002e4c424237365f36002e4c706372656c5f6869313635002e4c616e6f6e2e34313466363731613135666237623063306532636261396133343630323939342e3333002e4c706372656c5f6869313636002e4c616e6f6e2e34313466363731613135666237623063306532636261396133343630323939342e3334005f5a4e34636f726533666d7439466f726d6174746572323564656275675f7475706c655f6669656c64315f66696e6973683137683963326264643732306464613133376545005f5a4e34636f726533707472323864726f705f696e5f706c616365244c542424524624753634244754243137683536663832373834643464373061633345002e4c706372656c5f6869313637002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e343734005f5a4e37636b625f7374643130686967685f6c6576656c31396c6f61645f63656c6c5f6c6f636b5f686173683137686238376330343133623735373432633545005f5a4e37636b625f7374643130686967685f6c6576656c31346c6f61645f63656c6c5f646174613137686438663961623933373437336639633645002e4c706372656c5f6869313638002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e343330002e4c706372656c5f6869313730002e4c706372656c5f6869313639002e4c706372656c5f6869313731002e4c706372656c5f6869313732002e4c706372656c5f6869313733002e4c706372656c5f6869313735002e4c706372656c5f6869313734002e4c706372656c5f6869313736002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e3936002e4c706372656c5f6869313737002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e3234005f5a4e34636f7265336f70733866756e6374696f6e36466e4f6e63653963616c6c5f6f6e63653137683331326365396462383432326365623645005f5a4e34636f72653370747231303264726f705f696e5f706c616365244c542424524624636f72652e2e697465722e2e61646170746572732e2e636f706965642e2e436f70696564244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c542475382447542424475424244754243137683465633534623435323134663763393045002e4c43504938385f30005f5a4e34636f726533666d74336e756d33696d7037666d745f7536343137683238366534643532373433386334363745002e4c706372656c5f6869313738002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333234002e4c706372656c5f6869313739002e4c706372656c5f6869313830002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3233005f5a4e34636f726533666d7439466f726d617474657231327061645f696e74656772616c3137686238656639343965396131613633346545005f5a4e34636f726533666d7439466f726d617474657231327061645f696e74656772616c313277726974655f7072656669783137683834663538656430383761336264393345002e4c43504939315f30002e4c43504939315f31005f5a4e34636f726533666d7439466f726d6174746572337061643137683433336537613934646232626438653245002e4c706372656c5f6869313831002e4c706372656c5f6869313832005f5a4e34636f726533666d743577726974653137683537653362636463656237646630393145002e4c706372656c5f6869313833005f5a4e36305f244c5424636f72652e2e63656c6c2e2e426f72726f774572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137686163386261333334363731373261333845002e4c706372656c5f6869313834002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e313730005f5a4e36335f244c5424636f72652e2e63656c6c2e2e426f72726f774d75744572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683636336332373865383138373636393045002e4c706372656c5f6869313835002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e313731005f5a4e34636f726533666d74336e756d35335f244c5424696d706c2475323024636f72652e2e666d742e2e4c6f7765724865782475323024666f7224753230246936342447542433666d743137686632356530653835343735353364373145002e4c706372656c5f6869313836002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333232002e4c4350493130305f30002e4c4350493130305f31002e4c4350493130305f32005f5a4e36385f244c5424636f72652e2e666d742e2e6275696c646572732e2e50616441646170746572247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f7374723137686539366438303337316562386433343445002e4c706372656c5f6869313837002e4c706372656c5f6869313838002e4c706372656c5f6869313839002e4c706372656c5f6869313930005f5a4e34636f726533666d74355772697465313077726974655f636861723137686664666234386663643336373461323845005f5a4e34636f726533666d743557726974653977726974655f666d743137683364623431343565346436363932376245002e4c706372656c5f6869313931002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333237005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f7374723137683865303931326361326264646233386345005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e577269746524475424313077726974655f636861723137683239666437616639333939643762333645005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f666d743137683565373464633863623261616161323645002e4c706372656c5f6869313932005f5a4e34636f726533666d74386275696c64657273313044656275675475706c65356669656c643137686134393061356537663734366534656245002e4c706372656c5f6869313934002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e323933002e4c706372656c5f6869313935002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333030002e4c706372656c5f6869313933002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333031002e4c706372656c5f6869313936002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e323839002e4c706372656c5f6869313937002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e323932005f5a4e34636f726533666d74386275696c6465727338446562756753657435656e7472793137686531623638303262326163636539656445002e4c706372656c5f6869323031002e4c706372656c5f6869313939002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333033002e4c706372656c5f6869313938002e4c706372656c5f6869323030002e4c706372656c5f6869323033002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333032002e4c706372656c5f6869323032002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e313537005f5a4e34636f726533666d74336e756d35325f244c5424696d706c2475323024636f72652e2e666d742e2e55707065724865782475323024666f72247532302469382447542433666d743137683438643832613435336137306166353745002e4c706372656c5f6869323034005f5a4e34636f726533666d74336e756d35325f244c5424696d706c2475323024636f72652e2e666d742e2e4c6f7765724865782475323024666f72247532302469382447542433666d743137683039663834613031663936303437366145002e4c706372656c5f6869323035005f5a4e34325f244c54242452462454247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137686332303631326561373836393861653445002e4c706372656c5f6869323036002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333337005f5a4e36375f244c5424636f72652e2e61727261792e2e54727946726f6d536c6963654572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683532646436363362353834636335356645002e4c706372656c5f6869323037002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e353537002e4c706372656c5f6869323038002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e353333002e4c706372656c5f6869323130002e4c706372656c5f6869323039005f5a4e34636f726533666d74336e756d35335f244c5424696d706c2475323024636f72652e2e666d742e2e55707065724865782475323024666f7224753230246936342447542433666d743137683464336136353331313038303933376445002e4c706372656c5f6869323131005f5a4e35616c6c6f63377261775f7665633139526177566563244c542454244324412447542437726573657276653231646f5f726573657276655f616e645f68616e646c653137686332663335393562613638613033633645005f5a4e34325f244c54242452462454247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683035646461313430303562373034353645005f5a4e34325f244c54242452462454247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683431323134373832613466363464656645005f5a4e36355f244c5424616c6c6f632e2e7665632e2e566563244c5424542443244124475424247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137686464613861616433336135376363313045002e4c706372656c5f6869323132002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e323533002e4c706372656c5f6869323133002e4c706372656c5f6869323134002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333038005f5a4e35616c6c6f63337665633136566563244c54245424432441244754243131657874656e645f776974683137683935323361376565386561616133316645005f5a4e35616c6c6f63377261775f7665633139526177566563244c542454244324412447542437726573657276653231646f5f726573657276655f616e645f68616e646c653137686534386235666233366361343936633545005f5a4e35616c6c6f63377261775f766563313166696e6973685f67726f773137686465323762646133633136313431313345005f5a4e396d6f6c6563756c65323672656164657237726561645f61743137686436323832346538376630396538383045002e4c706372656c5f6869323234007374722e312e333135002e4c706372656c5f6869323137002e4c706372656c5f6869323138002e4c706372656c5f6869323135002e4c706372656c5f6869323136002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e31002e4c706372656c5f6869323233002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3136002e4c706372656c5f6869323235002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3139002e4c706372656c5f6869323139002e4c706372656c5f6869323230002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e36002e4c706372656c5f6869323231002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3132002e4c706372656c5f6869323232002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3134005f5a4e36315f244c54246d6f6c6563756c65322e2e7265616465722e2e4572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683238346238363235356264316239336545002e4c706372656c5f6869323236002e4c7377697463682e7461626c652e5f5a4e36315f244c54246d6f6c6563756c65322e2e7265616465722e2e4572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683238346238363235356264316239336545002e4c706372656c5f6869323237002e4c7377697463682e7461626c652e5f5a4e36315f244c54246d6f6c6563756c65322e2e7265616465722e2e4572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d7431376832383462383632353562643162393365452e343330002e4c706372656c5f6869323330002e4c706372656c5f6869323238002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e32002e4c706372656c5f6869323239002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e33002e4c706372656c5f6869323331002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3238005f5a4e396d6f6c6563756c65323672656164657236437572736f723133756e7061636b5f6e756d6265723137683635326430373132666263326536343145002e4c706372656c5f6869323332002e4c706372656c5f6869323333002e4c706372656c5f6869323334002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3331002e4c706372656c5f6869323335002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3335002e4c706372656c5f6869323432002e4c706372656c5f6869323336002e4c706372656c5f6869323337002e4c706372656c5f6869323431002e4c706372656c5f6869323338002e4c706372656c5f6869323339002e4c706372656c5f6869323430002e4c706372656c5f6869323433002e4c706372656c5f6869323434002e4c706372656c5f6869323435002e4c706372656c5f6869323436002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3430002e4c706372656c5f6869323437002e4c706372656c5f6869323438002e4c706372656c5f6869323439002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3538002e4c706372656c5f6869323530002e4c706372656c5f6869323531002e4c706372656c5f6869323532002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3634005f5a4e36395f244c5424616c6c6f632e2e7665632e2e566563244c54247538244754242475323024617324753230246d6f6c6563756c65322e2e7265616465722e2e526561642447542434726561643137683538323363346134366134643066373445002e4c706372656c5f6869323533002e4c706372656c5f6869323534002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3638005f5a4e34636f726533707472343664726f705f696e5f706c616365244c5424616c6c6f632e2e7665632e2e566563244c5424753824475424244754243137683139303635656264313265376238616645005f5a4e31387370617273655f6d65726b6c655f74726565346832353634483235363131706172656e745f706174683137683635373836666235326663646564306445005f5a4e37305f244c54247370617273655f6d65726b6c655f747265652e2e747265652e2e4272616e63684b6579247532302461732475323024636f72652e2e636d702e2e4f72642447542433636d703137683263653439633663323334323262346545005f5a4e39385f244c5424636b625f7374642e2e686967685f6c6576656c2e2e517565727949746572244c54244624475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137686231366136333531633137303061613745002e4c706372656c5f6869323535007374722e302e333530002e4c706372656c5f6869323537002e4c706372656c5f6869323536005f5a4e35616c6c6f6335626f7865643136426f78244c542454244324412447542431336e65775f756e696e69745f696e3137683834373362316265336534316438633545005f5a4e35616c6c6f6335626f7865643136426f78244c542454244324412447542431336e65775f756e696e69745f696e3137683761393538346163663734633633393245005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f646532313448616e646c65244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e4e6f6465526566244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4d75742443244b24432456244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e496e7465726e616c24475424244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e45646765244754243130696e736572745f6669743137686530613963663030393033343261333745005f5a4e35616c6c6f633131636f6c6c656374696f6e733562747265653673656172636839315f244c5424696d706c2475323024616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e4e6f6465526566244c5424426f72726f77547970652443244b24432456244324547970652447542424475424313466696e645f6b65795f696e6465783137683538623066623732343130626338653045005f5a4e35616c6c6f633131636f6c6c656374696f6e733562747265653672656d6f76653235395f244c5424696d706c2475323024616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e48616e646c65244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e4e6f6465526566244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4d75742443244b24432456244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4c65616624475424244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4b562447542424475424313472656d6f76655f6c6561665f6b763137683932356266653833663964336631323045005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b244324562447542432356d657267655f747261636b696e675f6368696c645f656467653137683565316662626261313330613939366445005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b2443245624475424313662756c6b5f737465616c5f72696768743137683134353762643930393139373763616445005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b2443245624475424313562756c6b5f737465616c5f6c6566743137686637323766663464373765333137663345005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b244324562447542438646f5f6d657267653137683764663761343032346566636539366545002e4c706372656c5f6869323538002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3731002e4c706372656c5f6869323539002e4c706372656c5f6869323631002e4c706372656c5f6869323630002e4c706372656c5f6869323632002e4c706372656c5f6869323634002e4c706372656c5f6869323633002e4c706372656c5f6869323635002e4c706372656c5f6869323636002e4c706372656c5f6869323638002e4c706372656c5f6869323637002e4c706372656c5f6869323639002e4c706372656c5f6869323730005f5a4e35616c6c6f6335626f7865643136426f78244c542454244324412447542431336e65775f756e696e69745f696e3137683865303536326639626532336432623745005f5a4e35616c6c6f6335626f7865643136426f78244c542454244324412447542431336e65775f756e696e69745f696e3137686630333839343435343838663831633145005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f646532313448616e646c65244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e4e6f6465526566244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4d75742443244b24432456244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e496e7465726e616c24475424244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e45646765244754243130696e736572745f6669743137683463363562306630323863663661333845005f5a4e35616c6c6f633131636f6c6c656374696f6e733562747265653673656172636839315f244c5424696d706c2475323024616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e4e6f6465526566244c5424426f72726f77547970652443244b24432456244324547970652447542424475424313466696e645f6b65795f696e6465783137686366633034636463626438393439336245005f5a4e35616c6c6f633131636f6c6c656374696f6e733562747265653672656d6f76653235395f244c5424696d706c2475323024616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e48616e646c65244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e4e6f6465526566244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4d75742443244b24432456244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4c65616624475424244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4b562447542424475424313472656d6f76655f6c6561665f6b763137686430343065343765356162316639336445005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f64653132354e6f6465526566244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4d75742443244b24432456244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4c6561664f72496e7465726e616c24475424313663686f6f73655f706172656e745f6b763137683662323932356361633530363230653245005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b244324562447542432356d657267655f747261636b696e675f6368696c645f656467653137683639343536653266653337656664353245005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b2443245624475424313662756c6b5f737465616c5f72696768743137683333636262626135643162656234643245005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b2443245624475424313562756c6b5f737465616c5f6c6566743137683565653138306237396130613266636245005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b244324562447542438646f5f6d657267653137683062356263386231666365346431343845002e4c706372656c5f6869323731002e4c706372656c5f6869323732002e4c706372656c5f6869323734002e4c706372656c5f6869323733002e4c706372656c5f6869323735002e4c706372656c5f6869323737002e4c706372656c5f6869323736002e4c706372656c5f6869323738002e4c706372656c5f6869323739002e4c706372656c5f6869323831002e4c706372656c5f6869323830002e4c706372656c5f6869323832002e4c706372656c5f6869323833005f5a4e34636f726535736c69636534736f727437726563757273653137686635623239333039636436333933336245005f5a4e34636f726535736c69636534736f72743235696e73657274696f6e5f736f72745f73686966745f6c6566743137683133346537316232363032303439623045005f5a4e34636f726535736c69636534736f72743134627265616b5f7061747465726e733137683038373030316334666161636539623445005f5a4e34636f726535736c69636534736f727432327061727469616c5f696e73657274696f6e5f736f72743137683664666664346137303338356239303045005f5a4e34636f726535736c69636534736f72743868656170736f72743137683739313663343261326535636431383945002e4c4350493136335f30005f5a4e35616c6c6f63377261775f7665633139526177566563244c54245424432441244754243136726573657276655f666f725f707573683137683266373139353338366332346364373445002e4c706372656c5f6869323834005f5a4e31387370617273655f6d65726b6c655f74726565356d65726765356d657267653137683733636631633763646362636630363645002e4c706372656c5f6869323837005f5a4e347574696c33736d7431316e65775f626c616b6532623137686530346638633332383130656566666645005f5a4e31387370617273655f6d65726b6c655f74726565356d6572676531304d6572676556616c756534686173683137686361663934316539633361336137646145002e4c706372656c5f6869323835002e4c706372656c5f6869323836005f5a4e31387370617273655f6d65726b6c655f74726565356d6572676531356d657267655f776974685f7a65726f3137686262316663663731613061663431616545002e4c706372656c5f6869323838002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3331002e4c4350493136395f30002e4c4350493136395f31002e4c4350493136395f32002e4c4350493136395f33002e4c706372656c5f6869323839002e4c706372656c5f6869323930002e4c706372656c5f6869323931002e4c706372656c5f6869323932002e4c706372656c5f6869323933005f5a4e34636f726535736c69636534736f72743236696e73657274696f6e5f736f72745f73686966745f72696768743137686537623533613633393836633665636245002e4c706372656c5f6869323934002e4c4350493137335f30005f5a4e35616c6c6f63377261775f7665633139526177566563244c54245424432441244754243136726573657276655f666f725f707573683137686331393061356231623136306436373545002e4c706372656c5f6869323935005f5a4e39385f244c5424636b625f7374642e2e686967685f6c6576656c2e2e517565727949746572244c54244624475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683639396362383835316633373032373345002e4c706372656c5f6869323936002e4c706372656c5f6869323937002e4c4a54493137355f30002e4c42423137355f31002e4c42423137355f32002e4c42423137355f33002e4c42423137355f34002e4c42423137355f35002e4c706372656c5f6869323938005f5a4e34636f726533707472373964726f705f696e5f706c616365244c5424636b625f7374616e64616c6f6e655f74797065732e2e67656e6572617465642e2e626c6f636b636861696e2e2e5363726970744275696c646572244754243137683230353465616461363664306463376345002e4c706372656c5f6869323939002e4c706372656c5f6869333030002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3437002e4c706372656c5f6869333032002e4c706372656c5f6869333031002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e313134002e4c706372656c5f6869333033002e4c706372656c5f6869333034002e4c706372656c5f6869333038002e4c706372656c5f6869333035002e4c706372656c5f6869333036002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3438002e4c706372656c5f6869333037002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e313139002e4c706372656c5f6869333132002e4c706372656c5f6869333039002e4c706372656c5f6869333130002e4c706372656c5f6869333131002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e313237002e4c706372656c5f6869333231002e4c706372656c5f6869333133002e4c706372656c5f6869333134002e4c706372656c5f6869333135002e4c706372656c5f6869333136002e4c706372656c5f6869333137002e4c706372656c5f6869333138002e4c706372656c5f6869333139002e4c706372656c5f6869333230002e4c706372656c5f6869333232005f5a4e347574696c3668656c70657232366765745f6d65746164615f646174615f62795f747970655f69643137683437383266333330623964363130353445002e4c706372656c5f6869333235002e4c706372656c5f6869333233002e4c706372656c5f6869333234002e4c706372656c5f6869333236002e4c706372656c5f6869333237002e4c706372656c5f6869333238002e4c706372656c5f6869333239002e4c706372656c5f6869333330002e4c706372656c5f6869333331002e4c706372656c5f6869333332002e4c706372656c5f6869333333002e4c706372656c5f6869333334002e4c706372656c5f6869333335002e4c706372656c5f6869333336002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3532002e4c706372656c5f6869333339002e4c706372656c5f6869333337002e4c706372656c5f6869333338002e4c706372656c5f6869333430002e4c706372656c5f6869333434002e4c706372656c5f6869333431007374722e32002e4c706372656c5f6869333432002e4c706372656c5f6869333433002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3439002e4c706372656c5f6869333439002e4c706372656c5f6869333538002e4c706372656c5f6869333539002e4c706372656c5f6869333639002e4c4a54493139315f30002e4c42423139315f333137002e4c42423139315f323530002e4c42423139315f323537002e4c42423139315f323631002e4c42423139315f323733002e4c42423139315f323739002e4c706372656c5f6869333436002e4c706372656c5f6869333438002e4c706372656c5f6869333631002e4c706372656c5f6869333632002e4c706372656c5f6869333633002e4c706372656c5f6869333735002e4c706372656c5f6869333733002e4c706372656c5f6869333630002e4c706372656c5f6869333634002e4c706372656c5f6869333635002e4c706372656c5f6869333636002e4c706372656c5f6869333531002e4c706372656c5f6869333532002e4c706372656c5f6869333435002e4c706372656c5f6869333437002e4c706372656c5f6869333637002e4c706372656c5f6869333638002e4c706372656c5f6869333530002e4c706372656c5f6869333536002e4c706372656c5f6869333537002e4c706372656c5f6869333533002e4c706372656c5f6869333534002e4c706372656c5f6869333535002e4c706372656c5f6869333731002e4c706372656c5f6869333732002e4c706372656c5f6869333730002e4c706372656c5f6869333736002e4c706372656c5f6869333734005f5a4e397374616b655f736d7431315f42554444595f484541503137686233373038373966306266356136656445005f5a4e397374616b655f736d7431375f46495845445f424c4f434b5f484541503137683263393037643763366462633565363545002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3134002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3237002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3732002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3733002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3734002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3735002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3736002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3737002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3738002e4c6c696e655f7461626c655f737461727430002e4c6c696e655f7461626c655f73746172743100626c616b6532622d7265662e63006c6f61643634002478007365637572655f7a65726f5f6d656d6f7279002478006d656d7365745f762e3000626c616b6532625f636f6d707265737300247800626c616b6532625f7570646174652e706172742e30002478002478002478002478002478002e4c3020002e4c3020002e4c3020002e4c3020002e4c3020002e4c3020002e4c3020002e4c3020002e4c3020002e4c34002e4c35002e4c3130002e4c3132002e4c3131002e4c3020002e4c3020002e4c3020002e4c3020002e4c3020002e4c3020002e4c3020002e4c3020002e4c3135002e4c3236002e4c3434002e4c3438002e4c3531002e4c3532006c69622e63002478002478002478002478002e4c32002e4c33002e4c3335002e4c3437002e4c3132002e4c3739002e4c3830002e4c3134002e4c3135002e4c3136002e4c3831002e4c3138002e4c3230002e4c3231002e4c3738002e4c3235002e4c3236002e4c3237002e4c3238002e4c3331002e4c3332002e4c3333002e4c3334002e4c3330002e4c3137002e4c3239002e4c3130002e4c313433002e4c313437002e4c313438002e4c313439002e4c323033002e4c313532002e4c323034002e4c313735002e4c313736002e4c313632002e4c323031002e4c313737002e4c313638002e4c313730002e4c313738002e4c313731002e4c313733002e4c313536002e4c313539002e4c313630002e4c313631002e4c313634002e4c323035002e4c313537002e4c313637002e4c313534005f5f636b625f7374645f6d61696e005f7374617274006d656d6d6f7665006d656d637079006d656d636d70006d656d73657400626c616b6532625f75706461746500626c616b6532625f66696e616c00626c616b6532625f696e69745f6b65795f776974685f706172616d00626c616b6532625f696e69745f706172616d000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000120000000000000060010100000000006001000000000000100d00000000000000000000000000001000000000000000000000000000000009000000010000001200000000000000700e010000000000700e000000000000400000000000000000000000000000000800000000000000080000000000000017000000010000000200000000000000b00e010000000000b00e000000000000c4170000000000000000000000000000080000000000000000000000000000002100000001000000060000000000000074360100000000007426000000000000be820100000000000000000000000000040000000000000000000000000000002700000001000000030000000000000038c902000000000038a9010000000000a8000000000000000000000000000000080000000000000000000000000000002e000000010000000300000000000000e0c9020000000000e0a9010000000000b8000000000000000000000000000000080000000000000000000000000000003400000001000000030000000000000098ca02000000000098aa010000000000080000000000000000000000000000000800000000000000000000000000000046000000080000000300000000000000a0ca020000000000a0aa01000000000000200800000000000000000000000000010000000000000000000000000000004b0000000100000000000000000000000000000000000000a0aa0100000000002802000000000000000000000000000001000000000000000000000000000000590000000100000000000000000000000000000000000000c8ac0100000000009c2600000000000000000000000000000100000000000000000000000000000065000000010000000000000000000000000000000000000064d3010000000000300200000000000000000000000000000100000000000000000000000000000074000000010000000000000000000000000000000000000094d5010000000000801300000000000000000000000000000100000000000000000000000000000082000000010000003000000000000000000000000000000014e901000000000012500000000000000000000000000000010000000000000001000000000000008d000000010000000000000000000000000000000000000026390200000000005d1c0000000000000000000000000000010000000000000000000000000000009d000000010000000000000000000000000000000000000083550200000000002400000000000000000000000000000001000000000000000000000000000000ad0000000300007000000000000000000000000000000000a7550200000000002b00000000000000000000000000000001000000000000000000000000000000bf0000000100000000000000000000000000000000000000d255020000000000041f000000000000000000000000000001000000000000000000000000000000cb0000000100000030000000000000000000000000000000d6740200000000002300000000000000000000000000000001000000000000000100000000000000d400000002000000000000000000000000000000000000000075020000000000c82d010000000000150000008d0c000008000000000000001800000000000000dc0000000300000000000000000000000000000000000000c8a2030000000000ee00000000000000000000000000000001000000000000000000000000000000e60000000300000000000000000000000000000000000000b6a3030000000000086c000000000000000000000000000001000000000000000000000000000000",
        "0x"
      ],
      "witnesses": [
        "0x55000000100000005500000055000000410000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0x"
      ]
    },
    "0xe6a4b80a06bbfbdb23456e6845b8ee87aa9644ad185c25295c919dbe6dbd8da0": {
      "version": "0x0",
      "cell_deps": [
        {
          "out_point": {
            "tx_hash": "0xf8de3bb47d055cdf460d93a2a6e1b05f7432f9777c8c474abf4eec1d4aee5d37",
            "index": "0x0"
          },
          "dep_type": "dep_group"
        }
      ],
      "header_deps": [],
      "inputs": [
        {
          "since": "0x0",
          "previous_output": {
            "tx_hash": "0x986220a6bafe37c3d7f8e2bb4dfbb7392188d142449cf38b098ba8b1a24009b6",
            "index": "0x1"
          }
        }
      ],
      "outputs": [
        {
          "capacity": "0x16d8d8708600",
          "lock": {
            "code_hash": "0x9bd7e06f3ecf4be0f2fcd2188b23f1b9fcc88e5d4b65a8637b17723bbda3cce8",
            "hash_type": "type",
            "args": "0x61a0d1fa2b4a4536a778659d5d87b88e82188b17"
          },
          "type": {
            "code_hash": "0x00000000000000000000000000000000000000000000000000545950455f4944",
            "hash_type": "type",
            "args": "0x3d8894c8397ff65858f87811ac394c0a0449f2a36ee21eae37ad597ed271cfa0"
          }
        },
        {
          "capacity": "0x149e0b67f2b00",
          "lock": {
            "code_hash": "0x9bd7e06f3ecf4be0f2fcd2188b23f1b9fcc88e5d4b65a8637b17723bbda3cce8",
            "hash_type": "type",
            "args": "0x61a0d1fa2b4a4536a778659d5d87b88e82188b17"
          },
          "type": null
        }
      ],
      "outputs_data": [
        "0x7f454c460201010000000000000000000200f30001000000cc340100000000004000000000000000c8cf0300000000000100000040003800050040001400120006000000040000004000000000000000400001000000000040000100000000001801000000000000180100000000000008000000000000000100000004000000000000000000000000000100000000000000010000000000cc24000000000000cc2400000000000000100000000000000100000005000000cc24000000000000cc34010000000000cc340100000000005c550100000000005c5501000000000000100000000000000100000006000000287a010000000000289a020000000000289a02000000000060010000000000006021080000000000001000000000000051e57464060000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000dc47010000000000fe4b010000000000a84f010000000000ac4f0100000000008c63010000000000aa9f010000000000bc9f010000000000ce9f010000000000e69f010000000000fc9f010000000000ee76020000000000988102000000000098810200000000009881020000000000c27802000000000098810200000000009881020000000000267b020000000000e27c020000000000327d020000000000617474656d707420746f206164642077697468206f766572666c6f770000000026a00100000000000000000000000000010000000000000042b301000000000046350100000000001800000000000000080000000000000036b601000000000026a001000000000001000000000000000100000000000000cab9010000000000617474656d707420746f206164642077697468206f766572666c6f770000000008c9bcf367e6096a3ba7ca8485ae67bb2bf894fe72f36e3cf1361d5f3af54fa5d182e6ad7f520e511f6c3e2b8c68059b6bbd41fbabd9831f79217e1319cde05b26a00100000000000000000000000000010000000000000042ab010000000000617474656d707420746f207368696674206c6566742077697468206f766572666c6f7700000000000000000000000000617474656d707420746f206d756c7469706c792077697468206f766572666c6f77000000000000000000000000000000617474656d707420746f2073756274726163742077697468206f766572666c6f77000000000000000000000000000000617474656d707420746f2073686966742072696768742077697468206f766572666c6f77000000000000000000000000617474656d707420746f206164642077697468206f766572666c6f776c6561662073697a65206d75737420626520616c69676e20746f20313620627974657300dc0301000000000023000000000000007265717569726573206d6f7265206d656d6f727920737061636520746f20696e697469616c697a65204275646479416c6c6f630000000000100401000000000033000000000000006f7574206f66206d656d6f72790000000000000000000000617474656d707420746f20646976696465206279207a65726f00000000000000617474656d707420746f206164642077697468206f766572666c6f7742797465735265616465725769746e65737341726773526561646572556e6b6e6f776e0026a001000000000008000000000000000800000000000000bab5010000000000456e636f64696e674f766572666c6f7776616c69646174654c656e6774684e6f74456e6f7567680026a001000000000008000000000000000800000000000000bab50100000000004974656d4d697373696e67496e6465784f75744f66426f756e6429426f72726f774572726f72426f72726f774d75744572726f725b000000aea201000000000018000000000000000800000000000000e0ab0100000000009cad01000000000050ae0100000000002020202052656164446174612c0a2c20280a282c0a5d30783030303130323033303430353036303730383039313031313132313331343135313631373138313932303231323232333234323532363237323832393330333133323333333433353336333733383339343034313432343334343435343634373438343935303531353235333534353535363537353835393630363136323633363436353636363736383639373037313732373337343735373637373738373938303831383238333834383538363837383838393930393139323933393439353936393739383939aea20100000000000800000000000000080000000000000088ae01000000000092ae01000000000048af0100000000002829000000000000aea2010000000000080000000000000008000000000000002cb301000000000054727946726f6d536c6963654572726f72636b622d64656661756c742d68617368616c726561647920626f72726f7765640000000000000026a00100000000000000000000000000010000000000000042ab010000000000616c7265616479206d757461626c7920626f72726f77656426a00100000000000000000000000000010000000000000030ab01000000000026a001000000000001000000000000000100000000000000cab90100000000000000000000000000617474656d707420746f206164642077697468206f766572666c6f77726561645f6174206069662073697a65203c20726561645f6c656e60726561645f6174206069662064732e63616368655f73697a65203e2064732e6d61785f63616368655f73697a6560726561645f617420606966206375722e6f6666736574203c2064732e73746172745f706f696e74207c7c202e2e2e60726561645f61742060696620726561645f706f696e74202b20726561645f6c656e203e2064732e63616368655f73697a656076616c69646174653a2073697a65203e206375722e736f757263652e746f74616c5f73697a65756e7061636b5f6e756d6265726765745f6974656d5f636f756e74636f6e766572745f746f5f753634636f6e766572745f746f5f753136636f6e766572745f746f5f7538636f6e7665727420746f205665633c75383e00000000007abf010000000000180000000000000008000000000000004ebe0100000000004669656c64436f756e744f75744f66426f756e64556e6b6e6f776e4974656d4f6666736574486561646572546f74616c53697a65436f6d6d6f6e617373657274696f6e206661696c65643a20696478203c204341504143495459000000000000000000000000000000000000000000000000000000000000000063616c6c656420604f7074696f6e3a3a756e77726170282960206f6e206120604e6f6e65602076616c7565000000617474656d707420746f206164642077697468206f766572666c6f7700000000617373657274696f6e206661696c65643a206f666673657420213d2030202626206f6666736574203c3d206c656e63616c6c65642060526573756c743a3a756e77726170282960206f6e20616e2060457272602076616c75650000000000000026a001000000000010000000000000000800000000000000949f01000000000046350100000000001800000000000000080000000000000036b601000000000026a00100000000000000000000000000010000000000000042b3010000000000617373657274696f6e206661696c65643a20656467652e686569676874203d3d2073656c662e686569676874202d2031617373657274696f6e206661696c65643a2073656c662e686569676874203e2030617373657274696f6e206661696c65643a207372632e6c656e2829203d3d206473742e6c656e2829617373657274696f6e206661696c65643a20656467652e686569676874203d3d2073656c662e6e6f64652e686569676874202d2031617373657274696f6e206661696c65643a20636f756e74203e2030617373657274696f6e206661696c65643a206f6c645f72696768745f6c656e202b20636f756e74203c3d204341504143495459617373657274696f6e206661696c65643a206f6c645f6c6566745f6c656e203e3d20636f756e74696e7465726e616c206572726f723a20656e746572656420756e726561636861626c6520636f6465617373657274696f6e206661696c65643a206f6c645f6c6566745f6c656e202b20636f756e74203c3d204341504143495459617373657274696f6e206661696c65643a206f6c645f72696768745f6c656e203e3d20636f756e74617373657274696f6e206661696c65643a206d6174636820747261636b5f656467655f696478207b5c6e202020204c6566744f7252696768743a3a4c6566742869647829203d3e20696478203c3d206f6c645f6c6566745f6c656e2c5c6e202020204c6566744f7252696768743a3a52696768742869647829203d3e20696478203c3d2072696768745f6c656e2c5c6e7d617373657274696f6e206661696c65643a206e65775f6c6566745f6c656e203c3d204341504143495459617373657274696f6e206661696c65643a20636865636b706f696e745f646174612e69735f6e6f6e652829617373657274696f6e206661696c65643a207374616b655f61745f646174612e69735f6e6f6e652829617373657274696f6e206661696c65643a2077697468647261775f61745f646174612e69735f6e6f6e65282906000000000000000900000000000000060000000000000006000000000000000b000000000000000a000000000000000a000000000000000400000000000000080000000000000004000000000000002c0901000000000023090100000000001d0901000000000017090100000000000c090100000000000209010000000000f808010000000000a805010000000000f804010000000000a4050100000000001000000000000000017a5200017801011b0c02001c00000018000000c62600006400000000420e2048810188028903920400000010000000380000000a27000010000000000000001c0000004c00000006270000ee00000000420e304a81018802890392049305002c0000006c000000d4270000d404000000420e80035a810188028903920493059406950796089709980a990b9a0c9b0d280000009c000000782c0000dc00000000420e6056810188028903920493059406950796089709980a990b0014000000c8000000282d00002c00000000420e104281010014000000e00000003c2d00002c00000000420e10428101002c000000f8000000502d00007a01000000420e900158810188028903920493059406950796089709980a990b9a0c00002c000000280100009a2e0000aa01000000420ea0015a810188028903920493059406950796089709980a990b9a0c9b0d2c0000005801000014300000c001000000420ed0015a810188028903920493059406950796089709980a990b9a0c9b0d2c00000088010000a43100008201000000420eb0015a810188028903920493059406950796089709980a990b9a0c9b0d2c000000b8010000f63200005002000000420ed0035a810188028903920493059406950796089709980a990b9a0c9b0d2c000000e801000016350000c600000000420e6058810188028903920493059406950796089709980a990b9a0c0000003000000018020000ac350000861e000000440ef00f74810188028903920493059406950796089709980a990b9a0c9b0d420ea010100000004c020000fe5300000a000000000e00001000000060020000f45300000a000000000e00001000000074020000ea5300000a000000000e00001000000088020000e05300000800000000000000100000009c020000d453000008000000000000001c000000b0020000c85300004e00000000420e304a810188028903920493050018000000d0020000f65300003000000000420e20468101880289030010000000ec0200000a54000008000000000000001000000000030000fe53000008000000000000001000000014030000f253000008000000000000001000000028030000e65300000800000000000000100000003c030000da5300000a000000000e00001400000050030000d05300000e00000000420e10428101001800000068030000c65300005800000000420e4044810188020000001800000084030000025400005800000000420e40448101880200000018000000a00300003e5400005800000000420e40448101880200000018000000bc0300007a5400005800000000420e40448101880200000018000000d8030000b65400005800000000420e40448101880200000018000000f4030000f25400005800000000420e40448101880200000018000000100400002e5500005800000000420e404481018802000000180000002c0400006a5500005800000000420e4044810188020000001400000048040000a65500005200000000420e40428101001800000060040000e05500005800000000420e404481018802000000140000007c0400001c5600005200000000420e40428101001800000094040000565600004e00000000420e30448101880200000018000000b0040000885600005800000000420e40448101880200000018000000cc040000c45600005800000000420e40448101880200000018000000e8040000005700008600000000420e30468101880289030018000000040500006a5700004c00000000420e30448101880200000018000000200500009a5700004e00000000420e304481018802000000180000003c050000cc5700009400000000420e6044810188020000001800000058050000445800009400000000420e6044810188020000001c00000074050000bc580000bc00000000420ee00348810188028903920400001c00000094050000585900009a00000000420e2048810188028903920400000020000000b4050000d2590000dc00000000440e304c8101880289039204930594060000002c000000d80500008a5a0000ee1a000000420ef0035a810188028903920493059406950796089709980a990b9a0c9b0d1c0000000806000048750000f000000000420e604881018802890392040000002c00000028060000187600001404000000420e80015a810188028903920493059406950796089709980a990b9a0c9b0d1000000058060000fc7900003c000000000e0000100000006c060000247a00000a000000000e000010000000800600001a7a00004c000000000e00001000000094060000527a00004c000000000e000010000000a80600008a7a0000f4000000000e00002c000000bc0600006a7b0000d403000000420eb00158810188028903920493059406950796089709980a990b9a0c00002c000000ec0600000e7f0000f203000000420ec0015a810188028903920493059406950796089709980a990b9a0c9b0d200000001c070000d0820000d600000000420e504e8101880289039204930594069507001800000040070000828300004a00000000420e104481018802000000140000005c070000b08300003200000000420e10428101001800000074070000ca8300006e00000000420e50468101880289030014000000900700001c8400003400000000420e104281010020000000a8070000388400006c00000000420e304c81018802890392049305940600000010000000cc0700008084000022000000000e000018000000e00700008e8400003a00000000420e20468101880289030020000000fc070000ac840000fc00000000420e404e81018802890392049305940695070010000000200800008485000042000000000e00002000000034080000b28500005000000000420e304c8101880289039204930594060000001c00000058080000de8500007400000000420e404881018802890392040000002000000078080000328600006400000000420e304c8101880289039204930594060000001c0000009c080000728600007a00000000420e2048810188028903920400000028000000bc080000cc8600009601000000420e900154810188028903920493059406950796089709980a000010000000e80800003688000072000000000e000014000000fc080000948800009200000000420e104281010010000000140900000e89000002000000000000001800000028090000fc8800007a00000000420e40448101880200000018000000440900005a8900008200000000420e4044810188020000002400000060090000c08900006001000000440ee008648101880289039204930594069507960897091000000088090000f88a000018000000000e0000100000009c090000fc8a0000040000000000000014000000b0090000ec8a00000e00000000420e104281010010000000c8090000e28a0000020000000000000014000000dc090000d08a00004201000000420e30428101002c000000f4090000fa8b0000e401000000420e705a810188028903920493059406950796089709980a990b9a0c9b0d001c000000240a0000ae8d00005600000000420e304a810188028903920493050024000000440a0000e48d00007803000000420e505281018802890392049305940695079608970900140000006c0a0000349100000e00000000420e104281010024000000840a00002a9100007e01000000420e80015081018802890392049305940695079608000010000000ac0a000080920000120000000000000010000000c00a00007e920000120000000000000014000000d40a00007c9200000e00000000420e104281010014000000ec0a0000729200000e00000000420e104281010014000000040b0000689200007000000000420e90014281012c0000001c0b0000c0920000bc01000000420e90015a810188028903920493059406950796089709980a990b9a0c9b0d140000004c0b00004c940000b400000000420e104281010014000000640b0000e89400003800000000420e4042810100100000007c0b0000089500000a0000000000000014000000900b0000fe940000b600000000420e104281010014000000a80b00009c9500003a00000000420e404281010020000000c00b0000be9500002001000000420ea0014e810188028903920493059406950720000000e40b0000ba9600000001000000420ea0014e81018802890392049305940695071c000000080c0000969700009800000000420e4048810188028903920400000014000000280c00000e9800000e00000000420e104281010014000000400c0000049800007200000000420e900142810114000000580c00005e9800007200000000420e900142810110000000700c0000b8980000160000000000000018000000840c0000ba980000a200000000420e40468101880289030014000000a00c0000409900007000000000420e90014281011c000000b80c0000989900005200000000420e304a810188028903920493050018000000d80c0000ca9900007c00000000420e5046810188028903001c000000f40c00002a9a00006200000000420e2048810188028903920400000010000000140d00006c9a0000360000000000000010000000280d00008e9a00003000000000000000180000003c0d0000aa9a00004c00000000420e10448101880200000020000000580d0000da9a00008600000000420e504c8101880289039204930594060000001c0000007c0d00003c9b00006800000000420e304a8101880289039204930500180000009c0d0000849b00007c00000000420e50468101880289030018000000b80d0000e49b00005200000000420e20468101880289030018000000d40d00001a9c00005600000000420e10448101880200000020000000f00d0000549c00008201000000420e504e81018802890392049305940695070010000000140e0000b29d0000280000000000000010000000280e0000c69d00006200000000420e10180000003c0e0000149e00006800000000420e30448101880200000014000000580e0000609e00003000000000420e104281010024000000700e0000789e00006601000000420e80015281018802890392049305940695079608970918000000980e0000b69f00006400000000420e30448101880200000018000000b40e0000fe9f00007800000000420e40468101880289030018000000d00e00005aa000007e00000000420e4046810188028903001c000000ec0e0000bca00000a200000000420e50488101880289039204000000180000000c0f00003ea100007a00000000420e20468101880289030020000000280f00009ca10000b200000000420e504c810188028903920493059406000000100000004c0f00002aa2000010000000000000001c000000600f000026a200008c00000000420e4048810188028903920400000010000000800f000092a200004a000000000000001c000000940f0000c8a200007200000000420e5048810188028903920400000010000000b40f00001aa30000c0000000000e000014000000c80f0000c6a300002400000000420e104281010014000000e00f0000d2a300002400000000420e10428101002c000000f80f0000dea300001401000000420e6058810188028903920493059406950796089709980a990b9a0c0000001000000028100000c2a400006c000000000000002c0000003c1000001aa500007e03000000420ed0035a810188028903920493059406950796089709980a990b9a0c9b0d100000006c10000068a8000068000000000e00002c00000080100000bca800000603000000420ec0015a810188028903920493059406950796089709980a990b9a0c9b0d2c000000b010000092ab0000e802000000420ec0015a810188028903920493059406950796089709980a990b9a0c9b0d2c000000e01000004aae0000d002000000420eb0015a810188028903920493059406950796089709980a990b9a0c9b0d2c00000010110000eab00000ae02000000420ea0015a810188028903920493059406950796089709980a990b9a0c9b0d140000004011000068b300002400000000420e1042810100140000005811000074b300002400000000420e1042810100280000007011000080b300002801000000420e6056810188028903920493059406950796089709980a990b00200000009c1100007cb400006800000000420e404e8101880289039204930594069507002c000000c0110000c0b400000403000000440ea00674810188028903920493059406950796089709980a990b9a0c9b0d10000000f011000094b7000066000000000e00002c00000004120000e6b70000c602000000440ef00474810188028903920493059406950796089709980a990b9a0c9b0d2c000000341200007cba00004602000000420eb0025a810188028903920493059406950796089709980a990b9a0c9b0d2c0000006412000092bc00008e02000000440ef00474810188028903920493059406950796089709980a990b9a0c9b0d2c00000094120000f0be00000202000000420e90025a810188028903920493059406950796089709980a990b9a0c9b0d2c000000c4120000c2c000003629000000440ec0046a810188028903920493059406950796089709980a990b9a0c9b0d18000000f4120000c8e900008c00000000420e504681018802890300200000001013000038ea0000cc01000000440ec0045881018802890392049305940600001c00000034130000e0eb0000f600000000440ec00454810188028903920493052000000054130000b6ec00005402000000440ee0045881018802890392049305940600002800000078130000e6ee00000604000000420ee00156810188028903920493059406950796089709980a990b2c000000a4130000c0f20000e809000000420ec00158810188028903920493059406950796089709980a990b9a0c000024000000d413000078fc00005001000000420e9001528101880289039204930594069507960897092c000000fc130000a0fd00000c03000000420ed0015a810188028903920493059406950796089709980a990b9a0c9b0d240000002c1400007c000100c803000000420ec001508101880289039204930594069507960800001c000000541400001c0401006a00000000420ea00348810188028903920400001800000074140000660401008c00000000420e5046810188028903001c00000090140000d60401007200000000420e5048810188028903920400000020000000b014000028050100ce02000000440e800658810188028903920493059406000018000000d4140000d20701003200000000420e10448101880200000028000000f0140000e80701001803000000420eb00256810188028903920493059406950796089709980a990b2c0000001c150000d40a01008c03000000420ef0025a810188028903920493059406950796089709980a990b9a0c9b0d2c0000004c150000300e01009003000000420e80035a810188028903920493059406950796089709980a990b9a0c9b0d2c0000007c150000901101004e04000000420e80035a810188028903920493059406950796089709980a990b9a0c9b0d20000000ac150000ae1501008601000000420e90014c81018802890392049305940600002c000000d0150000101701005602000000420ef0015a810188028903920493059406950796089709980a990b9a0c9b0d1800000000160000361901007801000000420ea001468101880289032c0000001c160000921a01005402000000420ef0015a810188028903920493059406950796089709980a990b9a0c9b0d2c0000004c160000b61c01006607000000440ea00674810188028903920493059406950796089709980a990b9a0c9b0d180000007c160000ec2301007400000000440eb0044c810188028903300000009816000044240100463a000000440ef00f74810188028903920493059406950796089709980a990b9a0c9b0d420e90110000000002452c00014697100000e780600f9308d00573000000011106ec22e826e44ae02a890869833589016385a5021766010003360653898db3b4c502998013048503086097800000e780402efd1413040405e5f80335890001cd03350900e2604264a2640269056117330000670003fde2604264a2640269056182800c6591c5086117330000670063fb8280797106f422f026ec4ae84ee4aa8508612dc903b9050183b98500630b09060144aa840de426846387090003340422fd19e39d09fe814419a80334052151c883598521850497300000e78080f68355a4212285e3f3b9fe850991cc8e09a29903b50922fd1491c403350522fd14edfc11c8814911a022857d1981442a84e31309fa39a8a2700274e2644269a269456182806387090003350522fd19e39d09fe8335052199c92e8497300000e78060f0833504212285e5f911a02a842285a2700274e2644269a269456117330000670043ee97300000e780c0ed17d5ffff130545349305b00297700000e780a0360000097186fea2faa6f6caf2ceeed2ead6e6dae25efe62fa66f66af26eee2a8a0061ae8a55c883348a008811a2852686d68697100000e780e0e80e75630605402e7b03b50a0083b50a014e7cee7d2af8aee003b58a0083b50a0203b68a0283bb8a012afc2ef032f463090b080359ab212d45138d0a026376a90c13851d006362a90213060003b385cd02da953305c5025a95b306b9413386c60297500100e780601603b50a0193050003b385bd02da9588e903b50a0088e103b58a0088e523bc750103350d0088f103358d001b04190088f5231d8b20a5a603b50a0183b50a00aae02ef803b58a0083b50a0203b68a0283bb8a012afc2ef032f497000000e780804b8355a5212d4663ffc5381b861500231dc520130600038666b385c5024276aa9594e9e27690e10276227794e523bc750190f198f52330aa0023340a00054511a622e405491545914c26e863eead006389ad000149994c63979d01814d954c21a0ee8c11a0e51d97000000e780a0448359ab212a8493c4fcffce94231d952013050003b385ac02da9588111306000397500100e78020c2314563f6a42c13851c00b385a9406397953013060003b305c502da953386c402228597500100e78080bf231d9b2108198c111306000397500100e78040beda8463130900a28452ec03d9a42113851d006362a90213060003b385cd02a6953305c5022695b306b9413386c60297500100e780c0ff03b50a0193050003130a0003b385bd02a69588e903b50a0088e103b58a0088e523bc750103350d0088f103358d00052988f5239d242188080c191306000397500100e78080b603350b216303051481449549a28a835c8b212a8b08018c081306000397500100e78040b4631b9c1e835dab212d4563e6ad1a0549114d63ee3c01668d638b3c01014919456395ac00814c154d19a0e51c194d97000000e780a0338359ab212a849344fdffce94231d9520b3054d03da9588111306000397500100e780a0ae314563faa418930b1d0033857941631e951813050003b385ab02da95130a00033386a402228597500100e780c0ab231dab2108198c111306000397500100e78080aa8359a42113851900b14563f4b9163386ad416316a616050c8e0bda9b93850b22930404220e06268597500100e78080a7014593153500a6958c6133363501239ca5203295b3b6a90093c61600758e23b8852065f288080c191306000397500100e78040a45a856313090022851001e685d68697000000e780201503350b21a28ae2849549e31505ec11a0014c97000000e7800024aa840355a5218145226623b0c42213890422139635004a961062b3b6a500231cb620b6953337b50013471700f98e23389620e5f2c26513851500626a23309a002334aa00639a850d83d9a4212945636c350d1b851900239da420130500033385a90226958c081306000397500100e780209a8509139539004a9500e123389420231c342111a810015a85e685d68697000000e780200a626a03350a0105052338aa00f6705674b6741679f669566ab66a166bf27b527cb27c127df26d19618280ad45268531a817d5ffff1305b5049305500315a017d5ffff1305550119a8b14597700000e7802077000017d5ffff1305f5ff9305800297700000e78060ec000017d5ffff1305a5e493050002edb717d5ffff1305b5fdf1bf17d5ffff130505f893050003c9bf17d5ffff130545e2e9bf1d7186eca2e8a6e4cae04efc52f856f45af05eec62e866e42a84835aa5213689b2892e8a93841500338bba4063e09a0213060003b305ca02a2953385c40222953306cb0297500100e78060ce938b1a00130500033305aa02229513060003ce8597500100e780c08793892a00130c042213052a00939c3400637c3501b3059c010e05629513163b0097500100e78020ca669c23302c01231d742163f434030e0a229a13058a22b305504109461461239c9620850423b88620b38695002105e397c6fee6604664a6640669e279427aa27a027be26b426ca26c25618280411106e413050022c14597300000e780c08f01c923380520231d0520a2604101828097300000e78040900000411106e413050028c14597300000e780008d01c923380520231d0520a2604101828097300000e780808d0000757106e522e1a6fccaf8cef4d2f0d6ecdae8dee4e2e066fc6af8aa8a0075035ca421330bbc002d45636b65112e8983bb8a0183d4ab2163ebb410338a2441239d4b21231d6421130d00033305a90322953306ac03a28597500100e78000ba930c1a00338594419305f9ff6318b50eb385ac03de95b309a50322854e8697400100e780c07203b50a0183b40a00330aaa035e9a3305a503aa940a8513060003a68597400100e7808070130600032685d28597500100e78060b4330534018a851306000397400100e780606e83b50a0203b50a03b9c541c9930404220e093385240113163c002106a68597500100e780e0b08e0ce69b93850b2226854a8697400100e780c06a0145050b8c601306150023b88520239ca520a1043285e317cbfe11a031e1aa600a64e6744679a679067ae66a466ba66b066ce27c427d4961828017d5ffff1305f5db930530031da017d5ffff130545de9305700221a817d5ffff1305b5d229a017d5ffff130535df9305800297700000e78080be0000357106ed22e926e54ae1cefcd2f8d6f4daf0deece2e8e6e4eae06efc2a89033b8501035cab212e8de2952d456363b5148339890203d5a9216364a515b30ca541231dbb20239d9921930bfdff930d00030335090103340900338abb03ae84b38a49013305b5032a940a8513060003a28597400100e780e05b130600032285d685a68a97500100e780a09f3305bc035a958a851306000397400100e780805993041c0033859a406392ab0e3385b4035a95ce85528697400100e780a057b305bd03ce953386bc034e8597500100e780409b8335090203350903adcd4dcd13840922139534005a951305052213193d00a2854a8697400100e780c053b305240113963c002106228597500100e780609763705c030e0c5a9c13058c220c61239c9520850423b865217d1d2105e3180dfe7d556382ac020145938b1c000c601306150023b83521239ca52021043285e397cbfe11a029e1ea604a64aa640a69e679467aa67a067be66b466ca66c066de27d0d61828017d5ffff130535c9930520030da017d5ffff130575cb11a817d5ffff130515b829a017d5ffff130595c49305800297700000e780e0a30000557186e5a2e126fd4af94ef552f156ed5ae95ee562e1e6fceaf8eef483bd850103dcad21628701c698750357a7216367d71632ec36f02af483ba850283dcaa21130b1c0033069b012d456360c516806188652ae488712ae883bb05010359a42132e0239dcd20130a0003b3844b03a294081813060003a68597400100e780c04093891b009385040313c5fbff330d250133064d03268597500100e780c08333054c036e950c181306000397400100e780a03d33054b036e9533864c03d68597400100e780603c93050422139539002e9593943b00a695c10513163d0097400100e780607f63f02903a294138584220c611386190023b88520239c35212105b289e317c9fe0315a4217d358545231da420226563f3a50413153b006e951305052293850a2213963c00210697400100e780a03502656372ac02850c0e0c6e9c13058c22da851061231cb62085052338b621fd1c2105e3980cfe626513341500568597200000e78020437d143375640182752e95a27523b0b501426690e588e9ae600e64ea744a79aa790a7aea6a4a6baa6b0a6ce67c467da67d6961828017d5ffff130595b19305100939a017d5ffff1305c5b99305a00297700000e780e0870000717106f522f126ed4ae94ee552e1d6fcdaf8def4e2f0e6eceae8eee4033a850183398502035baa2183dba92113041b0033067401ad4563ebc512833c05000c652ee4833d050103ddac2132e0231dca2013090003b38a2d03e69a080813060003d68597400100e780202693841d0093850a0313c5fdff330ca50133062c03568597400100e780206933052b0352950c081306000397400100e780002333052403529533862b03ce8597400100e780c02193850c22139534002e95939a3d00d695c10513163c0097400100e780c06463f0a403e69a13858a220c611386140023b89521239c95202105b284e317cdfe0395ac217d358545239dac20a26463f29504131534005295130505229385092213963b00210697400100e780001b02656371ab02850b0e0b529b13058b220c61239c8520050423b84521fd1b2105e3980bfe4e8597200000e78000296685a685aa700a74ea644a69aa690a6ae67a467ba67b067ce66c466da66d4d61828017d5ffff1305a5a19305a00297600000e780c06f0000457186e7a2e326ff4afb4ef752f356ef5aeb5ee762e3e6feeafaeef6ae8483bb050003ba05013289aa8983daab21130b000333046a035e940a8513060003a28597400100e7802010930504031345faff569533066503228597400100e7808053fd3a13950a03239d5b2183ba8400419195456372b51a2819de85568697800000e780a03a6a7505cd85456317b5068001080113068003a28597400100e780a00a6a65aa750355a52183d5a5212e950505b1456376b50408180c01014605a88001a80013068003a28597400100e780a0070675c6750355a52183d5a5212e950505b145637fb5020818ac000546d28697000000e78000bd89a80e65ae6599a0081a13068003a28597400100e780c003081a854597000000e78020a03665d66515a0050a081a13068003a28597400100e7808001081a854597000000e7804086766596752af82efcd2e0c27be27a03b60b21066a71c293841a00130b010c914d314c954c054d0354a62163e78d0a2819b285268697800000e780402b6a750dcd6318a509a81913068003da8597400100e78080fb526592750355a52183d5a5212e950505636c8503b3858c40a81997000000e780809691a8a81913068003da8597400100e78040f8526592750355a52183d5a5212e95050563728503081a13068003da8597400100e78000f6081a97000000e78020c92a86ae8409a8b3858c40a81997f0ffffe780a079014629fe29a001e405452300a9008a85130600034e8597400100e78040f223b8790323bc590323b04905be601e64fa745a79ba791a7afa6a5a6bba6b1a6cf67c567db67d796182801d7186eca2e8a6e4cae04efc52f856f45af05eec62e866e46ae0b289ae8a2a89938c0601130a0003854b130bf00f03dcaa21b3044c037d54568595cc130d050341055146e68597400100e780402d932505003335a000b305b040c98d938404fd05046a85e38b75fd13f5f50f631e65016396090089a06284638f09020e045694833a0422fd1965b701452334590123383901233c89002330a900e6604664a6640669e279427aa27a027be26b426ca26c026d256182802334590123380900233c89000545c9bf130101812334117e2330817e233c917c2338217d2334317d2330417d233c517b2338617b2334717b2330817b233c91792338a1792334b179797117560100130666570ce208e6081f1306004013040040814597400100e780c0d02330812405659b08a58105456215130715008c04081f01468146814701487300000039c1494413158403619545618330817e0334017e8334817d0339017d8339817c033a017c833a817b033b017b833b817a033c017a833c8179033d0179833d81781301017f8280833901241305104063e6a906854505444e8597700000e780e0f4aa8bae8a0c1f1306004097400100e78060d4938409c013850b402330912485659b88a5811317840305078c041306004081468147014873000000833501243335a000b3b5b4004d8d39c5e38c0af45e8597200000e780e0e0a9b74e85814597700000e78080eeaa8bae8a0c1f4e8697400100e78020ce114463ff89004545814597700000e78060ecaa842e8917c5ffff930575d889a003c51b0083c50b0003c62b0083c63b0022054d8d4206e206558e3364a60063998902214463f789084545814597700000e78040e8aa842e8917c5ffff930555d44546268597400100e78060c7054525a04545814597700000e780c0e5aa842e8917c5ffff9305d5d14546268597400100e780e0c401452328a13a233c813a2330313da8072334913c2338213dc545233cb13c0c6591c5086197200000e78000d34944e3860ae65e8597200000e78000d2b9bd03c55b0083c54b0003c66b0083c67b0022054d8d4206e206558e3364a6001335840093753400b335b0004d8d1dcd45454549814597700000e780a0dc2a84ae8417c5ffff9305b5c84546228597400100e780c0bb0d452328a13a281f233c813a2330913c2334213da5bf63ff89004545814597700000e780c0d8aa842e8917c5ffff9305d5c421b7135a24007d1a0d456377aa024545814597700000e78060d6aa842e8917c5ffff930575c24546268597400100e78080b511450d44c9a0631caa08114691445e85ce85a28697500000e780801913f63500f199b306b5002338a13a233cb13a2330d13c2334c13c2338913c88040c1f97500000e780e0f08804ce8597500000e780401803390124033401252338213b233c813a09452330a13c081f97500000e780a02921cd4545c549814597700000e780c0cc2a842e8917c5ffff9305d5b84546228597400100e780e0ab8d4441aa4545814597700000e78040caaa842e8917c5ffff930555b64546268597400100e78060a90d441145d28991b5e30c04100545e30ca41003360900833689005e85ce8597500000e780c00c99cd2a86ae86081fb285368697500000e78040118324013b15456399a4100945e303a40e03368900833609015e85ce8597500000e780400999cd2a86ae86081fb285368697500000e780c00d8324013b1545639da40c0d45e30da40a03360901833689015e85ce8597500000e780c00599cd2a86ae86081fb285368697500000e780400a8324013b15456391a40a0335812411c54a8597200000e78000ae938589ff0d456364b5006f10b00d938549ff6364b5006f10f00c03c59b0083c58b0003c6ab0083c6bb0022054d8d4206e206558eb366a60003c5db0083c5cb0003c6eb0003c7fb0022054d8d42066207598e3367a600081fde854e8697500000e780e0f5033a013c63020a080334013b5285814597700000e780c0b4aa842e89a285528697400100e78060948da0032a413b0334813b0339013c8339813c033b013d033c813d0335812419c50335012497200000e78080a22328913a232a413b233c813a2330213d2334313d2338613d0d45233c813d6387a40009456396a4008807c1b1281f75b9a80765b981440335813b19c50335013b97200000e780009e2944e38804ca0d45636445016f10700303c5140083c5040003c624008386340022054d8d4206e206558e518d85456315b50a081fa685528697500000e780c014033b013b0334013c2285814597700000e78040a72a8c2e8ada85228697400100e780e08619e06f10407e034b0c0063070a00628597200000e78040960335813b19c50335013b97200000e780209563070900268597200000e7804094054505496303ab000d49621513061500081f814597500000e780804c0345013b15c50335813b0e0597b5ffff938525572e950861054402850944f1bee30d09bc268597200000e780a08ff1b60315613b8315413b0356213b8346113b2312a10cc205d18d0334813b0335813c0356013d8334013caec12af9231cc10a638706360315410c8e45231aa1082ec91305610a0c19294697300100e780a07913550403231ea10813550402231da10813550401231ca108231b810813d504032312a10a13d504022311a10a13d504012310a10a231f9108081f0c09054697f00000e78020210334013b630404308304813b9305913b1305110d3d4697300100e7806073a2e52308910c8811ac0197200000e780c0c64e75930500026304b5006f10406b0e7583451500034605008346250003473500a205d18dc2066207d98ed58d034655008346450003476500834775002206558e4207e2075d8f598e0216d18daefd83459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2ee283451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2ee683459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5010345f5012206558e42076205598d518d02154d8d2aea081fac194a8697f00000e780e0cf0334013b6304041c8304813b9305913b130591243d4697300100e780005f2330812423049124081f8c040d4697700000e78020cd0339013b631409006f1040580305713c8305613c0346513c2307a136a205d18d2316b1360345213c8345113c0346313c8306413c22054d8d4206e206558e518d2324a1360345a13b8345913b0346b13b8346c13b22054d8d4206e2068345e13b558e518d0346d13ba2058346f13b0347013cd18d8304813bc2066207d98ed58d82154d8d2330a136228597700000e7806094130511128c163d4697300100e78080534aee23009112630b0b0e054549446317ab4813050002814597600000e780e0702a84ae89ac191306000297300100e7806050930500020546054a228597f00000e780e0a5aa8463870900228597100000e780205f13f5f40f130450046310454513050002814597600000e780006c2a84ae89ac191306000297300100e780804b930500020946228597f00000e78020a1aa8463870900228597100000e780605a13f5f40f8545130460046319b53e4a8597700000e780e0872e7511c50e7597100000e78000582e6597700000e780608663870a005e8597100000e780805601446ff04fea0d440db811443db039442db00344813b15b00344813b75a6081a2c0a97100000e780e07788042c0a97100000e780206c081f2c0a97100000e780e07003340124033601258334013b0337013ca802a285a68697d00000e780207e0335813b11c5268597100000e780804f0335812411c5228597100000e780804e88042c0a97100000e780c05b081f2c0a97100000e780806003340124033601258334013b0337013ca812a285a68697d00000e780c0780335813b11c5268597100000e780204a0335812411c5228597100000e780204928032c0a97100000e780e07188042c0a97100000e780a04a081f2c0a97100000e780604f03340124033601258334013b0337013c0813a285a68697d00000e780a0720335813b11c5268597100000e78000440335812411c5228597100000e7800043081fde854e8697500000e78020e48334013c95c08339013b2685814597600000e780404f2a8a2e89ce85268697300100e780e02e11a0014a0335813b19c50335013b97100000e780603e630f0a14081fd285268697500000e78000b88339013b8334013c2685814597600000e780804a2a842e8bce85268697300100e780202a23308124233461252338912488168c0497700000e780e0d50335813b19c50335013b97100000e780603863070900528597100000e7808037033501368335813603360137aae3aee7b2eba8020c091306000297300100e7800067012513046002631f0516081f0c09054697f00000e780e0ce8339013b6384090c0304813b9305913b1305111e3d4697300100e7802021ceef2300811e081f0c09094697f00000e780c0cb0335013baae845c50304813b9305913b1305911f3d4697300100e780001e4665aafb230c811ea80b97100000e780c05c9374f50f881b97100000e780e05b1375f50f130470026390a40e8804ac0b97100000e780006f081f8c1b97100000e780406e033601250335013c6315a6048335013b0335012497300100e780805a1339150015a84d447da80145814521a80545854509a80945894531a00344813b71a80d458d4597600000e78080f900000344813bbda801490335813b19c50335013b97100000e78040240335812419c50335012497100000e78020236306090413050002814597600000e78080302a8a2e8bac121306000297300100e7800010081f13060002d28597d00000e780807d0345013b3dc90344113b63070b00528597100000e780601e466597600000e780c04c4e8597600000e780204c1e6597600000e780804b5a6511c53a6597100000e780a01b727511c5527597100000e780c01a72694a8597600000e78000492e7511c50e7597100000e78020192e6597600000e78080476ff0afc50335813baae063070b00528597100000e7800017281e8c0397100000e78000722330013023380130281e97100000e780c063aae4630e051c814488162c1e268697100000e780c06a081f8c1697100000e780205c0335013cd1456304b5006f10e0000335013b83451501034605018346250103073501a205d18dc2066207d98ed58d2328b12483451500034605008346250003473500a205d18dc2066207d98ed58d034655008346450003476500834775002206558e4207e2075d8f598e0216d18d2330b12483459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f8336813b598e0216d18d2334b12489c697100000e78000078c045146880797300100e78040f588048c1697100000e7808039833501254145e399a5720335012403448500034b95000349a5008349b500034cc500834dd500834ce500034df50083450500aefc034a150083452500aef083453500aeec834545002ee583455500aef8834565002ee18335812403467500b2f489c597100000e780c0fe8504220b33658b004209e209b3e529014d8da20db3e58d01c20c620d33669d01d18d82154d8d220ae675b365ba0006764206e666e206558ed18d46762206aa66558e8a66c20626776207d98e558e0216d18d2338b13a233ca13a08060c1f97e0ffffe780800c0335013697600000e780a0262665e31795e283350131033681308336013003358133233cb1202338c1202334d12097600000e78000243e759e757e662338a1302334b1302330c130081f0c0697100000e78040270335013c93050002e315b5620335013b83459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18d233cb12483451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2338b12483459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2334b12483451500034605008346250003473500a205d18dc2066207d98ed58d034655008346450003476500834775002206558e4207e2075d8f8336813b598e0216d18d2330b12489c697100000e78040e1033581258335012503368124833601242334a13c2330b13c233cc13a2338d13a88168c0397100000e780203f8804866597f00000e780601428048c04101f941697f00000e780a01a058901e90335013097600000e780c00a21a82e840335013093f4f50f97600000e7808009e39d043e166593050002e318b54ad27703c5970183c5870103c6a70183c6b70122054d8d4206e206558e518d83c5d70103c6c70183c6e70103c7f701a205d18dc2066207d98ed58d82154d8d2334a13c03c5170183c5070103c6270183c6370122054d8d4206e206558e518d83c5570103c6470183c6670103c77701a205d18dc2066207d98ed58d82154d8d2330a13c03c5970083c5870003c6a70083c6b70022054d8d4206e206558e518d83c5d70003c6c70083c6e70003c7f700a205d18dc2066207d98ed58d82154d8d233ca13a03c5170083c5070003c6270083c6370022054d8d4206e206558e518d83c5570003c6470083c667003ee403c77700a205d18dc2066207d98ed58d82154d8d2338a13a88040c1f97e00000e78080c9033401246302047e0335012583358124130600053306c5022296233081222334b12232e8233cc1226305057e0665930525002eec33b5a5002af013050405aaf4880413068003a28597300100e780c0b2087c2ae1630d057803459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8d233ca1280345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8d2338a12803459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8d2334a1280345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8d2330a1280a652330a12a28642c1588e5286088e1081597100000e78020eb8275e3970518e265636cb566081f0c0597d00000e780203f0335013caaf863070566b007086a0c6610622330a12e233cb12c2338c12c4675233ca12a88050ce510e188162c1d97100000e78060eb081f8c1697100000e78000e08335013c4145e39da5180335013b034b850083499500834ca500034db5008344c500034cd5000344e5000349f50083450500aef0834d1500034a2500834535002efc834545002ee583455500aeec83456500aefc8335813b03467500b2e489c597100000e78060a5a20933e56901c20c620db3659d014d8d220cb3659c004204620933668900d18d821533e9a500a20d067533e5ad00420ae275e205b3e545014d8de665a2052a66d18d66764206a666e206558ed18d8215b3e4a500881697100000e78080ce1374f50f881697100000e78040d833e624018335013693461400558d3364a6002e8597600000e780e0cb631704549c1403c5170183c5070103c627018386370122054d8d4206e206558e518d232ca12e03c5970083c5870003c6a70083c6b70022054d8d4206e206558e518d83c5d70003c6c70083c6e70003c7f700a205d18dc2066207d98ed58d82154d8d2338a12e03c5170083c5070003c6270083c6370022054d8d4206e206558e518d83c5570003c6470083c6670003c77700a205d18dc2066207d98ed58d8215033d81204d8d2334a12e033b81213335a001833c0121b305a040b3f565012338a13a233c013a2330a13d2334913d2338a13c233c013c2330a13f2334913f2338b13e081f97600000e780204b69c5aa8413040501a8155146a28597300100e78060be012579fd0848906494600c0e88c9086088e1086488e5b6fc2330d13032e52334c130630b0d08281e1406ea85668697f0ffffe7806089033581333ded033501340336813483350135a30f0134630d06348e052e95033505229305f6ff89c90356a5210e06329503350522fd15edf98355a521fd15233ca1382330013a2334b13a081f2c0f1306f13597e0ffffe780c05e88160c1f1306000397200100e780e0710335013e8336013f8355a52163fcb6302a8605ae82fc02e5081f0c1597100000e780a0b48335013c41456392a56e0335013b0349850083499500034da5000344b5008344c500834cd500834de500034bf50083450500aee4034c1500834525002ef4034a350083454500aef0834555002efc83456500aeec8335813b0346750032f889c597000000e780007aa20933e52901420d6204b365a4014d8da20cb3e59c00c20d620b3366bb01d18d8215b3e4a500220c26653365ac00a275c205620ab365ba004d8de275a2050676d18d66664206c276e206558ed18d821533e4a500081597100000e78020a31375f50f85456315b502e675338585003336b500aa66b3859600b2956385d5002a6633b6c5006315065e014d014ba1a86675aa6563e395002285e6752e8d63e38500228daa65638395002a8d2a652a8b63639500268b667633358600aa66b38596403385a540018e6306d500aa65b3b5a50021a0e675b3b5c5009386f5ffb3f5a60033f5c6009814104b146718639c0790cb94e798e3233cb13a2338a13a28040c1f97d0ffffe780a07d33656d0163070514ba657a668816b415181397e00000e7802028081f8c16054697d00000e780e02e833c013c638b0c460334813bb00708620c66106a8334013b2330a1302334b1302338c13010170ce608e2233c9139081f8c16094697d00000e780202b8339013c638009440335813bac079061946598698335013b2330c1302334d1302338e130980614e710e3269db3369d00330664013696233c313363048600b3368600639b064ab345bd00318d4d8d631e053e280f97100000e780808c9374f50f281e97100000e780a08b1375f50f1304f007639ea43c08062c0f97100000e780408f081f2c1e97100000e780808e033601310335013c631da6008335013b0335013097300100e780408a1339150011a001490335813b19c50335013b97000000e78000570335813019c50335013097000000e780e055630c09364e8597600000e7800084668597600000e7806083467597600000e780c0820a6597600000e780208226752a84c265e31eb58c7da02330a136233401362338b136081f8c161306f13597e0ffffe780a02b25a88335813e0336052111ca835685210357a62185053285e3f7e6fe11a0ae86130500033385a60232958c161306000397200100e780403c0345f1357d1b233c6121e30a05ca638d0c3e03350d222334a120fd1c23389121233805206a8597000000e780404a41b903448124c5ac26740da026752338a12213041004f1a40344013b26752338a122c1a41304b0036da4426423388122081497d0ffffe780a044081397e00000e78080c993751500639405208335812003368121b336b00003370121b307d0407d8e2338d13a233c013a2330b13c2334e13c2338d13c233c013c2330b13e2334e13e2338c13e233c01321b5505012334013415cd931515002e957d15233ca13e081f97600000e780a0fc15c1aa8588041306000397200100e780a02d281e8c0497d0ffffe780e0510335813f79f588048c1b97000000e780c07003350125930500026313b52e0335012483459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18d233cb13683451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2338b13683459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2334b13683451500034605008346250003473500a205d18dc2066207d98ed58d034655008346450003476500834775002206558e4207e2075d8f83368124598e0216d18d2330b13689c697000000e780c02a03358137833501370336813683360136233ca1242338b1242334c1242330d12408068c0397100000e780e0918816866597e00000e780e05d281e8c169004140697e00000e7802064058911e9281e97d0ffffe780a02a29a81b54850039a02e84281e97d0ffffe78060291375f40f41e9280497d0ffffe7806028466597500000e78080511e6597500000e780e0505a6511c53a6597000000e7800021727511c5226597000000e780202072696fe09fc611456fe03ff90344013b05a00344013b01a8130400084e8597500000e780c04c668597500000e780204c26752338a122467597500000e780204b0a6597500000e780804a081497d0ffffe780e018280497d0ffffe780801f46656fe09ffc1145d2856fe03ff317a5ffff1305e55f9305b0028da017a5ffff1305e5e799a897400000e78040f1000017a5ffff1305856597a5ffff938625e89305b002100521a817a5ffff1305056497a5ffff9386a5ea9305b002100697400000e7800079000017a5ffff130525e329a017a5ffff130585e2f14597400000e780205c000041456fe05feb17a5ffff1305c55f97a5ffff938665e49305b002101f75bf17a5ffff1305455e97a5ffff9386e5e071b717a5ffff1305255d97a5ffff9386c5dfadbf17a5ffff1305055c97a5ffff9386a5dea5b717a5ffff130505679305100259bf97400000e78060e3000097400000e78080e4000097000000e78060ff0000173300006700e3bb173300006700a3f8797106f422f026ec4ae84ee43284ae892a89328597300000e780a0b9aa8405c163e38900a2892685ca854e8697200100e780c0f44a8597300000e780c0f42685a2700274e2644269a26945618280011106ec22e826e42a8497300000e78060b5aa8401c926858145228697200100e78000e42685e2604264a2640561828017030000670023f717030000670023f717030000670023f717030000670083fb97000000e78080f40000411106e497400000e78080d70000397106fc22f82a840a850d4697500000e780e05a02650dc14265a26502662af42ef032ec2c08228597600000e7802085e27042742161828017a5ffff1305454897a5ffff9386e5ce9305b002300897400000e780405d0000397106fc22f82a840a85114697500000e780605502650dc14265a26502662af42ef032ec2c08228597500000e780a07fe27042742161828017a5ffff1305c54297a5ffff938665c99305b002300897400000e780c0570000397106fc22f82a840a85154697500000e780e04f02650dc14265a26502662af42ef032ec2c08228597500000e780207ae27042742161828017a5ffff1305453d97a5ffff9386e5c39305b002300897400000e78040520000397106fc22f82a840a85194697500000e780604a02650dc14265a26502662af42ef032ec2c08228597500000e780a074e27042742161828017a5ffff1305c53797a5ffff938665be9305b002300897400000e780c04c0000397106fc22f82a840a851d4697500000e780e04402650dc14265a26502662af42ef032ec2c08228597500000e780206fe27042742161828017a5ffff1305453297a5ffff9386e5b89305b002300897400000e78040470000397106fc22f82a840a85214697500000e780603f02650dc14265a26502662af42ef032ec2c08228597500000e780a069e27042742161828017a5ffff1305c52c97a5ffff938665b39305b002300897400000e780c0410000397106fc22f82a840a85354697500000e780e03902650dc14265a26502662af42ef032ec2c08228597500000e7802064e27042742161828017a5ffff1305452797a5ffff9386e5ad9305b002300897400000e780403c0000397106fc22f82a840a85394697500000e780603402650dc14265a26502662af42ef032ec2c08228597500000e780a05ee27042742161828017a5ffff1305c52197a5ffff938665a89305b002300897400000e780c0360000397106fcaa852800014697500000e780002f226519cd6265c26522662af82ef432f0081097500000e7808051e2702161828017a5ffff1305a51c97a5ffff938645a39305b002101097400000e780a0310000397106fc22f82a840a85054697500000e780c02902650dc14265a26502662af42ef032ec2c08228597500000e7800054e27042742161828017a5ffff1305251797a5ffff9386c59d9305b002300897400000e780202c0000397106fcaa852800094697500000e7806024226519cd6265c26522662af82ef432f0081097500000e780603fe2702161828017a5ffff1305051297a5ffff9386a5989305b002101097400000e78000270000797106f422f02a840a85194697500000e780201f026519c94265a265026608e80ce410e0a27002744561828017a5ffff1305450d97a5ffff9386e5939305b0021306f10197400000e78020220000397106fc22f82a840a85094697500000e780401a02650dc14265a26502662af42ef032ec2c08228597500000e7808044e27042742161828017a5ffff1305a50797a5ffff9386458e9305b002300897400000e780a01c0000397106fc22f82a840a85014697500000e780c01402650dc14265a26502662af42ef032ec2c08228597500000e780003fe27042742161828017a5ffff1305250297a5ffff9386c5889305b002300897400000e78020170000797106f422f026ec0c6911466394c500814491a0006110600865050610e031c21306450022e06360a6040d4532e46371b504f1152ee80a8597500000e780e0fc0a8597500000e780e008aa84228597500000e78080db2685a2700274e264456182800000000017a5ffff130505f229a017a5ffff130565f19305b00297400000e780c0f30000797106f422f02a840a8597500000e7800007026519c94265a265026608e80ce410e0a27002744561828017a5ffff130525f59795ffff9386c57b9305b0021306f10197400000e780000a0000797106f422f02a840a85014697500000e7802002026519c94265a265026608e80ce410e0a27002744561828017a5ffff130545f09795ffff9386e5769305b0021306f10197400000e780200500001d7186eca2e82a842818054697500000e78040fd627539c12665866562762aec2ee832e408102c0097500000e780e011027529c14275a2750276aae4aee032fc2c18228597500000e780c0252265e6604664256117530000670023c917a5ffff130565e89795ffff9386056f9305b002101021a817a5ffff1305e5e69795ffff9386856d9305b002301897400000e780e0fb00001d7186eca2e82a842818094697500000e78000f4627539c12665866562762aec2ee832e408102c0097500000e780a008027529c14275a2750276aae4aee032fc2c18228597500000e780801c2265e66046642561175300006700e3bf17a5ffff130525df9795ffff9386c5659305b002101021a817a5ffff1305a5dd9795ffff938645649305b002301897400000e780a0f20000057186efa2eba6e7cae3ae842a899385050828001306800f97100100e780807a9385040408021306000497100100e780607903b4841739cc038504001b05f5fb1375f50f1335050c9335140493c515004d8d39e52800a68597000000e780400613060008018e88022295814597100100e780606888020c02228697100100e780607428008c021306000897000000e780c00c39a02800a68597000000e78040022c001306800f4a8597100100e7808071fe605e64be641e693d618280011106ec22e826e44ae02e892a84130505041306800b814597100100e780e0611795ffff9305055913060004228597100100e780606d13053900a14522868346e5ff0347d5ff8347f5ff83440500a206d98ec207e204c58f0347150083442500dd8e834735000217a214458fc217830445005d8f1c62d98ee214c58ebd8e14e2fd1521062105c5fd0345090068f4e2604264a26402690561828069ce797106f422f026ec4ae84ee452e03284ae842a89687193050008b389a54063f6c9082330090e130a09065295a6854e8697200100e78060a80335090493050508033689042330b904133505f81345150032952334a9044a85d28597000000e78000083304344113051008ce94636fa402930900080335090493050508033689042330b904133505f81345150032952334a9044a85a68597000000e7804004130404f893840408e3e789fc0335090e4a9513050506a685228697200100e780e09f0335090e22952330a90ea2700274e2644269a269026a45618280417186f7a2f3a6efcaebcee7d2e356ff5afb5ef762f366ef6aeb6ee72e892a842801130600082401814597100100e78060490d0941458345e9ff0346d9ff8346f9ff03470900a205d18dc206620703461900d98e03472900d58d0216834639002217598e03074900c216558ed18d6217d98d8ce07d15a104210955fd280213060004a28597100100e780a0502c603064833204053267b2772a65aae89736010083b4e6b2033884053e972a97a58db98d9734010083b424b293d605028215d58d338e9500b346fe004a652ae193d78601a216dd8e2a973303d700b345b30013d70501c215b3e8e500469eb345de0093d6f50386055267d274ea67bee4173501000335e5adb3ebd50026973e97318d398d9735010083b525ad135605020215518daa95ad8c8a7636f813d68401a214d18c3386e600330996003345a900935605014215b36cd500338abc0033459a009355f5030605f26672772a769734010083b404a9b369b500ba96b296328c32f433c59200358d9734010083b4e4a79357050202155d8daa94258fca752eec935787012217d98fae96b382f60033c5a200935605014215b36dd500ee94a58f13d5f703860792761666ea75aefc17370100033707a433eba700b296ae963345e800358d17370100033727a39355050202154d8d2a97398e8e67bef0935586012216d18dbe96b383b60033c5a300135605014215518d2a97b98dae6a13d6f5038605d18d56934e933345a300135605020215498eb29433c53401ce69935685012215c98e338569004ee8b30ed50033c6ce00935706014216336df600b3009d0033c6d0006e6f9356f6030606b36fd6007a99fae033032b01b347130193d407028217c58f3e97b34467010e75aaf493d88401a21433e61401b3086500b298b3c7f80093d40701c21733e39700330be3003346cb002e75aaf81357f6030606b364e600aa92ae9233c69201135706020216598e329eb345be004e7913d78501a2154d8fb30559004af03388e5003346c800935206014216b36256003386c201318fee751355f7030607336ea700ae93ae86aeecde9333c5b301935d050202153365b501b30c4501b3cd7c01926793d58d01a21db3e5bd00be933e873efcb38db30033c5ad00935305014215336a750033059a01a98d93d7f5038605dd8db69eae9eb3c76e0093d607028217dd8e3696b18d93d78501a215dd8db387ee01b38eb700b3c6de0093d70601c216b3e3f6003383c300b345b30013d6f5038605b3ecc500e298fe98b3c5120113d605028215d18d2e953346f501935686012216d18e56e4338658013696b18d93d70501c215b3e8f500b382a80033c5d2009355f50306054d8d4e982698b3450a0193d605028215cd8eb690b3c5900093d78501a215cd8fb3050701b38ff500b3c6df0093d40601c21633e89600c290b3c6f00093d7f6038606d58fca9df29db3c6ad0193d406028216d58c338f6401b346cf0113d78601a216558fe676ee96338ae600b3449a0093d50401c214c58d2e9f3347ef009354f7030607d98c8a66b69eaa9eb3c5be0013d705028215d98d33871500398d935685012215c98e467b33856e01b30ed500b3c5be0013d50501c215b3eba500338deb00b346dd0013d5f6038606b3e0a600466c62963e96334576009355050202154d8d2a9fb345ff0093d68501a215d58d266e7296b309b60033c5a900935605014215558d2a9fb345bf0093d6f5038605b3edd5002676b29fa69fb3c51f0193d605028215cd8e3693b345930093d48501a215cd8c8675fe95b3839500b3c6d30093d70601c216d58f3e93b346930093d4f6038606b3e8960062673a9a669ab3460a0193d406028216c58eb692b3c4920193d58401a214c58d4279b3044901b38fb400b3c6df0093d40601c21633ea9600b3045a00a58d93d6f5038605d58db29eae9e33c5ae00935605020215c98eb382660033c5b200935585012215c98d33855e01b30cb500b3c6dc0013d50601c216b3eea600f69233c5b2009355f50306053363b50033063b010696b18f13d5070282175d8d3388a400b345180093d68501a215d58d62962e96318d935605014215b360d50006983345b8009355f50306054d8dba93ee93b3457a0093d605028215cd8eb387a601b3c5b70113d78501a215b3e4e500b385c301338a9500b346da0013d70601c216b3e3e6009e97bd8c93d6f4038604c58ee275ae9fc69fb3c47f0113d704028214458f3a9fb3441f0193d58401a214c58d827bde9fae9f33c7ef00935407014217458f3a9fb345bf0093d4f503860533ec95008665ae9caa9c33c7ec00935407020217458fba973d8d935485012215c98ce669338599012695298f935807014217336b1701b30cfb0033c79c009357f7030607b36df700ca8a4a96b305d60033c7be009357070202175d8fb307ef00bd8e93d48601a216c58e66762e96338dc6003346ed00135706014216b36ee600338efe00b346de0013d7f603860633efe6000676329a629a33471a00935407020217458fba92b3c5820193d48501a215cd8c8a68b3854801338a95003347ea00935707014217336cf700e292b3c7920093d4f7038607b3e097004267ba9f9a9fb3c77f0093d407028217c58f3e98b344680093d68401a214c58e2279ca9fb69fb3c7ff0093d50701c217dd8db3870501bd8e93d4f6038606c58e329536953346d501935406020216458e33085600b346d80093d48601a216c58e3a953695298e935406014216336396001a983346d8009356f6030606b362d600569d6e9d3346ac01935606020216d18eb69733c6b701135786012216598e3387a801b30ac700b3c6da0093d40601c216b3e39600b38df30033c6cd009356f6030606558e5e9a7a9ab3c5450193d605028215cd8eb3889601b3c5e80193d78501a215cd8fc675d295338ab700b346da0093d40601c21633ef9600fa98b3c7f80093d4f7038607c58fa675ae9f869fb3c66f0193d406028216d58cb38ec401b3c61e0093d58601a216d58db3863f01b38fb600b3c49f0093d60401c214c58eb69eb3c5be0093d4f5038605c58da66b5e953307c500b98e93d406028216c58eb69833c6c800935486012216458e66753a953295a98e93d40601c21633ec9600b30c1c0133c6cc009356f6030606336ed600e26833871a013e9733466700935606020216558e3303d601b346f30093d78601a216dd8e866a5697330dd7003346cd00135706014216598e3293b346d30013d7f6038606b3e0e600ca894a9a2e9ab3467a0013d706028216d98e3698b345b80013d78501a215d98dc66433079a00b38ee500b3c6de0093d70601c216dd8e3698b345b80093d7f5038605b3e3f5006279ca9f969fb3c5ef0193d705028215cd8fbe9db3c55d0013d78501a2154d8f226bb305fb01338fe500b347ff0093d50701c217dd8dae9d33c7ed009357f70306075d8fc2673e953a95298e9357060202165d8e32983347e8009357870122175d8f2695b307e5003d8e135506014216b362a60016983345e8001356f5030605518d2ae8469d729d33c5a601135605020215498eb29d33c5cd01935685012215c98e06756a95330dd5003346cd00135706014216b36fe600338ebf013346de009356f6030606d18ede9e869eb3c5d50113d605028215d18db388950133c61800135786012216598e33873e01b30dc700b3c5bd0093d40501c215b3ee9500f698b3c5c80013d6f50386054d8e569f1e9fb3458f0193d405028215cd8c2693b345730013d58501a2154d8db3052f01b383a500b3c4930093d50401c214c58db3846500258d1357f5030605498f6665aa97b697bd8d13d5050282154d8daa98b3c5d80093d68501a215d58d8a66be96b380b60033c5a000935705014215336af500b30b1a0133c5bb009355f50306053363b50026794a9d329d33c5a201935505020215c98db388b40033c5c800135685012215498e467c33058d01330fc500b345bf0093d70501c215cd8fbe98b3c5c80013d6f5038605b3e2c500667dea9dba9db3c5fd0113d605028215d18d2e983346e800135786012216518f33866d01da89b30ce600b3c5bc0093d40501c215c58d2e983347e8009354f7030607b36f9700c27dee934265aa9333c7d301935407020217d98cb38ac40133c7aa00135587012217598d027e33077e00b30ea700b3c49e0013d60401c214d18c33865401318d9356f5030605558da666b690aa90b3c6f00093d706028216dd8eb38a060133c5aa009357850122155d8db3878001aa97bd8e13d70601c21633e8e600c29a33c5aa009356f5030605b363d5006a9f1a9f33c5e501935505020215c98d2e9633456600935685012215c98e06657a95330dd500b345bd0013d70501c21533e3e500330fc300b345df0013d6f5038605d18d4665aa9c969c33c69401935606020216558eb29bb3c65b0013d78601a216558fb3862c013309d7003346c900935406014216336b9600da9b33c6eb001357f6030606598ece9efe9e33c74e01935407020217d98ca69833c7f801935687012217d98e3387be01330cd700b3449c0013d70401c214458fb3041701a58e13d5f6038606c98e2275aa97ae973d8f135507020217598db30f7501b3c5bf0013d78501a215d98df297338ab7003345aa00135705014215b362e500969f33c5bf008e689355f5030605b369b500469d329d33450d019355050202154d8db30e950033c6ce00ca7d135786012216598eb384ad01338dc4003345ad00135705014215498fba9e33c6ce00926c9357f6030606b36bf60066993699334669009357060202165d8eb29ab3c6da0093d78601a216dd8ee667ca97338ed7003346ce00135506014216518daa9a33c6da009356f60306063369d6008a652e9c1e9c33468b01935606020216d18e369f33467f004e68935786012216d18f33060c01338bc700b346db0013d60601c216558eb306e601b58fae7493d5f7038607dd8dd294ae94258f9357070202175d8f330f5701b3c5e50193d78501a215cd8fb385b401338cb70033478701935407014217336a9700529f33c7e701ca679354f703060733639700ea97ce973d8d135705020215598db303d500b3c6790013d78601a216558fb3869701b30cd70033459501935705014215b369f500ce93334577006e779357f50306055d8d72975e97398e9357060202165d8eb29fb3c7fb014e7e93d48701a217c58f7297338de7003346a601135706014216b36ae600d69f33c6f7012a779357f60306065d8e5a974a97b3c5e20093d705028215cd8fbe9eb345d901ee6693d48501a215cd8cb305d700b382b400b3c7570093d60701c217dd8eb69e33c7d401aa679354f7030607d98ce297aa97bd8e13d706028216d98eb69f3345f501135785012215598dc697330cf500b3c6860113d70601c21633e9e6004ae3ca9f3345f501ea761357f5030605b36be500e696b2963345da00135705020215598d330ad501334646018a7e135786012216598ef696b30dd6003345b501935605014215558d2a9a334646019356f6030606336bd600429d269d33c6a901935606020216558e329fb3c6e401ea6493d58601a216d58db3069d00b38cd50033469601935406014216458e329fb3c5e501ae6493d7f5038605b3e9f500a6929a92b3c55a0093d705028215cd8fbe93b34573008e7493d68501a215cd8eb3859200b38ab600b3c7570193d50701c217dd8db3877500bd8e13d7f6038606d98e629e369e3345c501135705020215598db302e501b3c6560013d78601a216d98e269e338cc60133458501135705014215b363e5009e9233c556009356f5030605336fd5007af6ee98de9833451601135605020215518d3303f50033c66b00ee76135786012216598ec696b30bd60033457501935605014215336ed5007293334566002e769356f5030605558d66965a96b18d93d605028215d58db386f5013347db00ca67935487012217d98c3e96338bc400b3c5650113d60501c215b3efc500fe96b58c93d5f4038604b3ecb400d69ece9eb345d90113d605028215d18d2e9a33c64901935486012216d18c33860e01b38ac400b3c5550113d60501c215d18d2e9a33c64401ca741357f6030606598ee294aa94a58d13d705028215d98dae96358d2a679357850122155d8d2697330de500b3c5a50113d70501c215b3eee50076e3b388de0033451501126c9356f50306053369d500e29be69b33c57301935605020215c98eb383460133c57c002a77935785012215c98f3385eb00338aa700b3c6460113d70601c216558fba93b3c677002e6893d7f6038606b3ebf600429b329bb3466e0193d706028216d58fbe9233465600ea75935686012216558eb306bb00330bd600b3c7670113d50701c2175d8daa92334656006a6e9357f6030606b369f600f29afa9a33c65f01935706020216d18f3e9333466f00ee66935486012216d18c3386da002696b18f93d60701c217dd8e3693b3c7640093d4f7038607c58fea95be952d8f935407020217d98ca69233c75700935787012217d98fe295b38ab700b3c4540193d50401c214b3efb400fe92b3c5570093d7f503ee74860533eff5007af6d294ca94258d935505020215c98d2e9333456900ce67135785012215498f3385f400330ca700b3c5850193d70501c21533eaf5005293b34567000e7793d7f5038605cd8f5a975e97b98e93d506028216d58dae98b3c61b018a7413d58601a216558d2697b304e500a58d93d60501c21533e9d500ca9833451501aa659356f5030605558db295ce9533c6be00935606020216558eb293b3c6790013d78601a216d98ec2953388b60033460601135706014216598eb293b3c676002e7793d5f6038606d58d56973e97398e935606020216558eb298b3c6170193d78601a216d58fb306c701b389d70033463601135706014216b36ee60076e3f69833c617014e779357f6030606336bf60062972a9733c6ef00935706020216d18fbe93334575008e6f135685012215518d3306f701330cc500b3c7870113d70701c2175d8fba93334575004a6e9357f5030605b36af500f294ae9433459a009357050202155d8daa92b3c555002a7a13d68501a215d18dd294b38c950033459501135605014215336dc500ea92b3c555006e6693d6f5038605b3ebd50032987a98b345090193d605028215cd8eb3846600b3459f004a7393d78501a215cd8fb30568003389b700b3c6260193d50601c216d58dae94a58f93d6f7038607dd8e4e963696318f9357070202175d8f33085700b3c60601ea6713d58601a216558d3e96b30dc5003347b701135607014217b369c7004e98334505011356f5032e670605336fc5007af662975a973345ed00135605020215518db302950033465b009357860122165d8e5297330be60033456501135705014215336ae500d292334556001356f5030605518de69fd69fb3c5f50113d605028215d18d3387150133c6ea00ea74935786012216d18f33869f00b38fc700b3c5f50193d40501c215b3e895004697b98f93d5f7038607dd8d4a9e5e9eb3c7ce0193d407028217c58fbe93b3c47b0013d68401a214458e7293b30e6600b3c7d70193d40701c217c58fbe933346760092649356f6030606558eee94aa94a58f93d607028217dd8e3383e600334565000e779357850122155d8d2697b30be500b3c6760193d70601c21633eef60072e3729333456500ce669357f50306053369f500da96ae9633c5d900935705020215c98fbe9333c57500ee75935485012215c98c3385b600338ba400b3c7670193d50701c217dd8dae93b3c674008a7a93d7f6038606b3e9f600d69fb29fb346fa0193d706028216dd8e369833460601ae77935486012216458efe97330cf600b3c6860193d40601c216c58e369833460601ce741355f6030606336aa600a69efa9e33c5d801135605020215518daa9233465f002a67935486012216458eba9e330fd6013345e5019357050142155d8daa92334656009357f60306065d8e5e973297b98d93d705028215dd8d2e9833460601ca67935486012216d18c3306f700b38cc400b3c5950113d70501c215b3efe5007e98b3c5040113d7f503ea678605b3eee50076f6da97ca97bd8e93d506028216cd8eb3885600b345190113d78501a2154d8fb3855701330bb700b3c6660193d70601c216b3eaf600d69833471701aa779354f7030607458fe297ce973d8d935405020215458d2a93b3c46900ca7693d58401a214c58dbe96b38bd500334575019356050142153369d5004a9333c56500ea759356f5030605c98efa95d2953345be00935405020215c98ca69333457a008e67135685012215498e3385f500330ca600b3c4840193d50401c214c58db38775003d8eae629354f6030606458e969cba9cb3c5950193d405028215c58db3836500334777004e63935487012217458fb3846c00330d9700b3c5a50113d50501c21533efa500fa9333457700ee6c9355f5030605b369b500669b369b33c56f019355050202154d8daa97bd8e8e7513d78601a216d98eda95338bb60033456501135705014215498f330ef70033c5c601ae769357f5030605336af500de96b29633c5da009357050202155d8d2a9833460601ce7f935786012216d18f3386f601b38bc70033457501935605014215558d2a98b3c50701ee7793d6f5038605b3ead5003e9c769cb345890193d605028215d58dae98b3c41e01926613d68401a214458eb304dc0033099600b3c5250193d40501c215c58dae98334616019354f6030606458eea97b2973d8f935407020217458f3a9833460601935486012216458ee697330cf60033478701935407014217b36e97007698334606011357f6030606aa74598e7ae332f6da94ce94258d135605020215518d3306150133c7c900935787012217d98f33875400b389e70033453501935405014215b36895004696b2ea3d8e1355f6030606b367a6005e93529333c565009355050202154d8daa93b3457a0013d68501a215d18d3306d3003383c50033456500935605014215b362d500969333c575009355f5030605b366b500ca9fd69f3345ff01935505020215c98d2e9e33c5ca01ea74135685012215498e33859f00330fa600b3c5e50193d40501c215cd8c269eb345c6014a6613d5f5038605c98d62963e96b18c13d504028214458daa93b3c77700ae7413d78701a2175d8f26963a9632e6318d135605014215518d2ae31e95aaee398d1356f5032a670605518d2afa4e97369733c5ee00135605020215518d2a9e33c6c601ea669357860122165d8eba96b29636ea358d935605014215558daaf67295aaf2318d1356f5038e760605518d2afe9a96ae9633c5d800135605020215518d2a98b3c505010e6613d78501a215d98d36962e9632ee318d135605014215518daafa4295aae62d8d9355f50306054d8daae23275ca75aa95fa9533c6b200d666135706020216598eb296358d0a779357850122155d8dba95aa952ef2b18d13d60501c215d18daefeb695aeea2d8d9355f5030605c98da8022ef6a1451060833605fc1861358e398e10e0fd1521052104f5f5be701e74fe645e69be691e6afa7a5a7bba7b1a7cfa6c5a6dba6d7d6182801d7186eca2e8a6e4cae02e89aa840a8513060004814597000100e780c09be8749305000263e9a50aa86855e5e870ac603386a500b46403c7040fb335b600b0e0b695ace419c3fd55acecfd5513061008ace86378c50813060008138404066309c500098e2295814597000100e780a0962685a28597e0ffffe780e04921459305310026861462a38ed5fe13d78600238fe5fe13d70601a38fe5fe13d786012380e50013d70602a380e50013d786022381e50013d70603a381e500e1922382d5007d152106a1055dfdf0748a854a8597000100e780209de6604664a6640669256182809305000897300000e78000800000197186fca2f8a6f4caf0ceecd2e8d6e4dae05efc62f866f46af06eec906103bc8500329c636fcc34aa8988699376f50093b616003337a000f98e6380063a814a89466368d5008d462a87850a0581e3ede6fe83cb85013285d68597000000e780a03b6365ac322a8d1305000463f5aa323305ac4133555501814c89456368b5008d452a86850c0581e3edc5fe938d2c0063ea9d316145b3b5ad02639a0530b384ad02ea9463eaa43113893c006a847d19268a630d0902630c0d24233044015285639b0b00130600105285814597000100e78060810860610408e1c10408e5e3f844fd1785ffff1305a589a5ac4ee0638b0d2e014b13098d0093891c005a85ee8597000000e780a03563030d201d05935435002330490163990b0052858145268697f00000e780207cd29463e24425638669016109050b268ad1b7094963e72d0593098d02330a904105442285ee8597000000e780c0301d05135b350023b0990063990b00268581455a8697f00000e780807733856401636195200504b3058a00e109aa84e39325fd11a02685d68597000000e7806028636fac2463860d262a8b938bfdff2a84638b0b161385edff9305f00363eda520854c5a846ae86ee463080d14aa843395ac00331d55013309a401636589186145b38da402c265ae9d3385ab022e9593098500130a0501636f2c0d03b50d000c612300b40013d68503a303c40013d605032303c40013d68502a302c40013d605022302c40013d68501a301c40013d605012301c400a181a300b40093558503a307b400935505032307b40093558502a306b400935505022306b40093558501a305b400935505012305b40093558500a304b4002304a4000c6180e500e15a85d6852686a28697000000e780c022058915ed5a85d6855e86a28697000000e780802183b5090013563500b295838605001d893395ac00c98e2380d50083350a00b29503860500518d2380a5004a846a99e37489f249a82685a26597000000e780c0185a85d6852686a28697000000e780801c83b58d0013563500b295038605001d893395ac00518d2380a50081cc1385f4ffa68b426de31c0dea97200000e78000e10000426da26d63638c0a33058c40826523b0650123b4850188e923bca50123b0b50323b45503e6704674a6740679e669466aa66a066be27b427ca27c027de26d096182801775ffff13052562f14597200000e780c0bf00001775ffff1305e560f5b71775ffff13054560cdb71775ffff1305a55fe1bf1775ffff13050559ada81775ffff1305655b93054002c9b71775ffff1305855d5dbf1775ffff1305e553a1a81775ffff1305455c4db71775ffff1305a55591a01775ffff1305054f9305300271b71775ffff1305255e29a85285d68597000000e780c002637bac001775ffff1305056197000000e780400500001775ffff130565519305100289bf01cd1306000463f0c5027d153355b50005053315b50082801775ffff1305054f9305100239a01775ffff130525519305400297200000e780a0b1000097100000e780c040000063efa5006382a5021345f5ffaa951305000463f2a50205453315b50082801775ffff1305454a29a01775ffff1305a5499305100239a01775ffff1305c5429305300297200000e78040ac000063e0a6041307f003636cc7001307000463fde500898e33d5c6003355b50082801775ffff1305654829a01775ffff1305c5479305400297200000e78040a800001775ffff1305e552b545f5b790659461137806fc3698636bd80c98699355660063e3e500ba8594e2094694e6b68763ebc508fd1593d8860393d2060313d3860293d3060213de860193de060113df8600b68736863e879387070463efe7062380c70013578603a383e700135706032383e70013578602a382e700135706022382e70013578601a381e700135706012381e7002182a380c7002384d700a387170123875700a386670023867700a385c7012385d701a384e70190621ce6fd159ce23e86c9f99385070463e7f50214e1233405010ce914ed82801775ffff1305e53bf14597200000e780809900001775ffff1305a53af5b71775ffff1305053acdb7717106f522f126ed4ae94ee552e1d6fcdaf8def4e2f0e6eceae82a841305000497150100138a65a863718504171501009304a5a78860631e05348864fd558ce063130512c870cc6cd068d464aae4aee032fc36f80a850c1897000000e780209c054588e413850401c5a803350a04631b053203358a04fd552330ba041ded03350a0883358a0703360a07aae02efc32f80a850c1897000000e78080e705452334aa040265a2654266e2662338aa04233cba042330ca062334da0603398a0663000902033509000c6110650ce20c6510610ce6130b0a04630825032a8991a403390a0603358a056373a902130509046368252983350a042330aa0685052330ba046315092209a823340a0619ac03350a0405052330aa0403350a00631e052803358a00fd552330ba001ded03350a0a83358a0903360a0983368a08aae4aee032fc36f80a850c1897000000e780408d05452334aa0013050a018a851306000397f00000e780c02683398a031305f003636335210545814c3315350163788500850c63840c1c0605e36c85fe83350a0363e3bc00e68503358a020146e146b386dc02aa96138406fdb385bc406389c516630d051c147803b9060061047d16e307d9fe033509008335890088e1033589008335090088e5047017150100130b058d03350b0183358b03934af6ffe69a5686ca8697000000e78000cd93553500a695038605001d89854b3395ab00518d2380a50063f85c11130c000417150100130be588138afaff63778a1333954b01b3143501ca9463e72413033d840203350b0183358b035686ca8697000000e780a0c793553500ea95038605001d893395ab00518d2380a500833a840003350b0183358b035286ca8697000000e780c0c493553500d695038605001d893395ab00518d2380a50008600c612380b40013d68503a383c40013d605032383c40013d68502a382c40013d605022382c40013d68501a381c40013d605012381c400a181a380b40093558503a387b400935505032387b40093558502a386b400935505022386b40093558501a385b400935505012385b40093558500a384b4002384a4000c6184e504e12114d28ae3e54cf119a00149528b03350b0005052330ab004a85aa700a74ea644a69aa690a6ae67a467ba67b067ce66c466d4d6182801775ffff1305e50421a81775ffff130545f89305300231a01775ffff13056503f14597100000e780006100001775ffff130525f6f9bf1775ffff13058501cdb797100000e780007b00001775ffff1305d5339775ffff9386c5f115a01775ffff1305b5329775ffff9386a5f009a81775ffff130595319775ffff938685efc1450a8697100000e78000760000317106fd22f926f54af14eed52e956e55ae1defce2f8e6f4eaf0eeec97050100938c656b83b50c04639d05382a8903b58c04fd5523b0bc041de9170501001304856948602c7c3078aae4aee032fc28002c1897000000e78060ae054528e42265c2656266827628e82cec30f034f403b50c0583b58c053335a9001345f5ffb335b9006d8d51c5170501001305c5642c75638e052090612300c90093568603a303d900935606032303d90093568602a302d900935606022302d90093568601a301d900935606012301d9002182a300c90013d68503a307c90013d605032307c90013d68502a306c90013d605022306c90013d68501a305c90013d605012305c90013d68500a304c9002304b900906165a203b50c0483b50c00050523b0ac04639b052a03b58c00fd5523b0bc0015ed170501001304455a48704c6c50685464aae8aee4b2e036fc28002c1897f0ffffe780c04f054508e4130504012c001306000397f00000e78060e983ba0c03638f0a2283b98c02138afaff13848902854463809a04638b0922033b040003b50c0183b58c032686ca8697000000e780609593553500da9583c505001d8933d5a50005898504610469d5f91463e6440139a263030a108144930a0004268b63e49a00130b000483bb8c0303bc0c0161453385a4024e9513048502054d03b50c0183b58c032686ca8697000000e780808f638e091a833504fe13563500b2950386050093767500b316dd0093c6f6ff758e2380c500937515003306b040833604fe13661600329513563500369603460600937675003356d600058a51e2630b9b1263fe5b1333159500331575016295636e85131061146590e21065146190e691c12a89833d040003b50c0183b58c0385042686ca8697000000e780c08693553500ee95038605001d893315ad001345f5ff718d2380a5006104e3129af4d28405a023302901930585064a862334260123b02501930c050451a8638a090e814461453385a4024e9508610c612300b90013d68503a303c90013d605032303c90013d68502a302c90013d605022302c90013d68501a301c90013d605012301c900a181a300b90093558503a307b900935505032307b90093558502a306b900935505022306b90093558501a305b900935505012305b90093558500a304b9002304a9000c6123b425012330250103b50c00050523b0ac00ea704a74aa740a79ea694a6aaa6a0a6be67b467ca67c067de66d296182801775ffff130545b829a01775ffff1305a5b79305300231a01775ffff1305c5c2f14597100000e780602000001775ffff130585bb93051002edb797100000e780c03a00001775ffff130595f39775ffff938685b109a81775ffff130575f29775ffff938665b0c145300097100000e780e03600005d7186e4a2e026fc4af84ef452f056ec83ba050263800a0a2e8a2a898065b35954034e8597000000e780200b83340a002ae02ee402e863e335078145636e54031396350032950d466370560983c6140003c70400a206d98e03c7240083c7340033045441d6944207e2075d8fd98e14e185052105e37a54fd2ee8226502662338b9002334a9002330c900a6600664e2744279a279027ae26a616182800a8581454e8697000000e780e007c2650265e37954f9d9b71775ffff1305c5bce54597100000e780600f00001145d68597200000e780e0970000411106e422e02a840dc51355c4030de993351500131534008e0511c597d0ffffe78080c1aa8599e597d0ffffe780c0c20000a1452e85a285a26002644101828097d0ffffe780e0c10000411106e497000000e780e002fd55fe1585056315b500a2604101828011e597d0ffffe78060bf000097d0ffffe78020be00005d7186e4a2e026fc2e966374b600014591a82a8408659314150063639600b284914563e39500914493d5c40393b51500139634008e0501c914600e0536f0a14636f42af811a002f42800141097200000e78040b9a265426591e508e004e47d557e150505a6600664e27461618280411106e4054697000000e780c0f8fd55fe1585056315b500a2604101828011e597d0ffffe78040b5000097d0ffffe78000b40000797106f422f026ec4ae84ee452e06365d7046366e604aa89b304d7403389d5002685814597200000e78020be2a842e8aca85268697f00000e780c09d23b0890023b4490123b89900a2700274e2644269a269026a456182803685ba8519a03a85b28597100000e780407f000063e8c60063e9d500b385c640329582803285b68511a0368597100000e780207d0000011106ec22e826e42a8410690865ae846319a6002285b28597000000e78060f210680860931536002e9504e1050610e8e2604264a26405618280397106fc22f826f44af04eec52e856e4114a32892a84637d46032d45ad4a814597200000e780e0b1aa84ae891775ffff9305459d2d46268597f00000e7800091054508c0233444012338240104ecb1a803c5150003c6050083c6250083c535002205518dc206e205d58db3e4a500b9c09104638424052d45ad4a814597200000e78020ac2a8aae891775ffff930585972d46528597f00000e780408b2320040004e423382401233c4401233034032334540331a0114a631d4901154508c0e2704274a2740279e269426aa26a216182802d45ad4a814597200000e78080a6aa84ae891775ffff9305e5912d46268597f00000e780a08523200400a9b71061833805011c65210605483e8763ee17019307f7ff10e11ce5637d1801833686ff0c622106e3f3d5fe333517011345150082800545854597100000e780a0650000797106f422f026ec4ae84ee452e02e89aa8413050002130a0002814597200000e780409e2a84ae8913060002ca8597e00000e780c07d80e023b4340123b84401a2700274e2644269a269026a45618280397106fc22f826f44af0b2841106636996042e892a843285814597200000e78060992ae02ee402e826ce10100a856c0897100000e780a07e330699000a85ca8597100000e780a07d4265a265026608e80ce410e0e2704274a2740279216182801765ffff1305657ff14597100000e78000d00000797106f422f026ec4ae84ee452e08d4663f3c604aa899304c6ff138945002685814597200000e780a0912a842e8aca85268697e00000e780407123b0890023b4490123b89900a2700274e2644269a269026a456182801145b28597100000e78020530000011106ec22e826e44ae02a841305000285451309000297c0ffffe780207d29c9aa8413060002814597e00000e780c05e04e0233424012338240111458545914497c0ffffe780807a05c5a301050023010500a30005002300050008ec04f004f423080402e2604264a26402690561828097c0ffffe78080790000757106e522e1a6fccaf8cef4d2f0d6ecdae8dee4e2e003bb050193040b0163e86415938b140063890b142e8a83ba8502b3895b0163e779152a894e85814597200000e78000822ae42ee802ec0d4597000000e780c0ae2af02ef402f899c1814501a8081097000000e78000bcc27502758e052e95c1450ce1c27585052ef822756398a500081097000000e780e0b9c275027c13953500629504e19384150026f82275639aa4000810a68597000000e780a0b7c274027c1394340033058c00233075014ede900028006c1897100000e780e05fa2797d556384a402930b0104210462850c61930485002ede28006c185e8697100000e780805d611426857df063870900628597c0ffffe780206783350a0013040a0333866501280097100000e780e05a13061a032800a28597100000e780e05983358a0133865501280097100000e780c0586265c26522662338a9002334b9002330c900aa600a64e6744679a679067ae66a466ba66b066c496182801765ffff1305655911a81765ffff1305c55829a01765ffff13052558f14597100000e780c0a800000d476371c7069306c6ff637ad704930686ff0d476375d70403c8550003c7450083c7650083c6750022083367e800c207e206dd8ed98e03c8950083c8850083c2a50083c7b500220833671801c202e207b3e757005d8f170300006700c3a61145b68519a01145b28597100000e780002b0000411106e410610e069766ffff9386c61e369610620286907588711c6e9765ffff938535593d4635a8907588711c6e9765ffff938565572d462da021052ae01765ffff930765531765ffff1307e5533d463da0907588711c6e9765ffff938545502146a2604101828721052ae01765ffff9307854c1765ffff1307854c1d468a862e85be8597100000e780a018a260410182808280397106fc22f83287ae862a8402f002ec02e802e4130500022af405659b0815822c108d472800894201460148730000006309550285456308b502914515e522751306000289456361a602130514002c001306000297e00000e78080372300040009a8854511a081450ce408e805452300a400e270427421618280397106fc22f83287ae862a8402f002ec02e802e4130500022af405659b0815822c109547280089420146014873000000630b55028545630cb502914515e922751306000289456365a602130524002c001306000297e00000e780e02f01458545a300b40009a80145a300040029a081450ce408e805452300a400e270427421618280130101ba233c1144233881442334914423302145233c3143233841432334514323306143233c7141b289ae8b2a8408081306004093040040814597e00000e780801c2338914005659b08c58293050141080889440146de864e8781470148730000006301950885456300b508914535ed03390141130500406372250b8545054b4a8597100000e78040442a8aae8a0c081306004097e00000e780c023930209c013050a402338514085659b88c58293050141130600408944de864e87814701487300000063019508630e6507114b25ed03350141094b63e8a2062330440123345401b1a8854511a081450ce408e8233004008330814503340145833481440339014483398143033a0143833a8142033b0142833b81411301014682804a85814597100000e780603aaa84ae890c084a8697e00000e780001a04e0233434012338240145bf014b2334640108e823300400e3810afa528597c0ffffe780802851bf9308d0057d558145014681460147814701487300000001a0086101a0411106e497c0ffffe780a01a00008280797106f42e8813564500130f7002130710279766ffff938e662f6363e608130f70021307610217f600008338a67939661b03068f05669b03b6479302c0f937e6f5051b0ef60faa86333515032d813b066502b307d600139607034992330676029355160141821376e67fbb855502be95769683471600c615c19103460600a30ff7fef69583c7150083c50500711f230fc7fea300f7002300b7007117e365defa130630066370a60493150503c99105661b06b647b385c502c5811306c0f93b86c502329546154191791f7695034615000345050093061100fa96a380c6002380a6002e85a945637cb5009305ffff130611002e961b0505032300a60005a006059305efff7695034615000345050093061100ae96a380c6002380a60093061100ae96130770020d8f1765ffff9305855e4285014697000000e780e000a27045618280597186f4a2f0a6eccae8cee4d2e056fc5af85ef462f066ec6ae86ee4aa8403654503ba893689328aae8b937c1500b70a110063840c00930ab00293754500ce9c89e5814b8c6085e5a1a08145630e0a005286de86038706008506132707fc134717007d16ba957df6ae9c8c6095c103bd840063ffac01218925ed83c58403054633059d41634cb60af9e1aa8c2e85c9a0807084742285a6855686de86528797000000e7806014054b0dc15a85a6700674e6644669a669066ae27a427ba27b027ce26c426da26d656182809c6c2285ca854e86a6700674e6644669a669066ae27a427ba27b027ce26c426da26d6561828780581305000383c584032ee003bc040283bd840288d8054b238c64036285ee855686de86528797000000e780e00c51f5228a33049d4105047d1451c803b60d02930500036285029665d985bf09466398c50093051500058193dc150011a0814c03bc040203bd84028458130415007d1409c803360d026285a68502966dd9054b2dbf37051100054be389a4f26285ea855686de86528797000000e780e00511fd83368d016285ca854e86829619f5b30990417d5a7d59338529016309450303360d026285a6850296050975d50da083b68d016285ca854e868296e31005ee014b23a844030265238ca402c1bd6689333b9901e1b5797106f422f026ec4ae84ee49b070600370811003a89b6842e84aa896389070114704e85b2858296aa85054591ed81cc1c6c4e85a6854a86a2700274e2644269a269456182870145a2700274e2644269a269456182805d7186e4a2e026fc4af84ef452f056ec5ae85ee483320500146933e7d2003289ae896304072a638706101c6d8146338e29018507370311009308f00d1308000f4e8601a893051600918eae962e866303640efd17adc7630fc60d8305060013f4f50fe3d105fe834516009374f40113f7f50363fa8802834526001a0793f5f503b363b7006367040383453600f614ad909a0393f5f50333e4b300458c630c64089305460055b79305260013946400598c61bf93053600b20433e4930071b7630bc6078305060063d3050493f5f50f1307000e63ede5021307000f63e9e50203471600834726001377f70393f7f70303463600f615ad9132079a075d8f1376f603598ed18d370611006386c50285c263fd2601b385d90083850500130600fc63d7c500814591e539a0e39d26ffce8599c13689ae89638b021803388500930500026372b902814e63060916ca85ce86038606008506132606fc13461600fd15b29efdf581aa13877900619b3386e940b308c90093f678008145630d3701ce87038407008507132404fc934414000506a6957df6014691ce93f788ffba9783840700850793a404fc93c41400fd162696fdf693d6380097f7000083b7872997f4000083b28429b714001092048504939804018508b30eb6001da013173e001a97b386c34113763e00b3f45500a181b3f55500a695b3851503c191ae9e2deaddcab6833a839305000c368e63e4b600130e000c9375ce0f139435001a94dddd81451a8745df146393c4f6ff9d8099821067c58efd8eb6959346f6ff9d82046b1982558e7d8e93c6f4ff9d829980c58e046ffd8e3696b29513c6f4ff1d829980458e7d8e13070702b295e31d87fabdb7630803029305000c63e4b3009303000c814593f633008e06106021041347f6ff1d831982598e7d8ee116b295f5f611a0814533f65500a181b3f55500b295b3851503c191ae9e63fc0e01834685030546b305d8416345d60285ce814a25a80c7508719c6dce854a86a6600664e2744279a279027ae26a426ba26b6161828709466398c600138615008581935a160019a0ae8a8145033b0502833b85020459138415007d1409c803b60b025a85a68502966dd9054a81a037051100054a638ca40283b68b015a85ce854a86829605e533095041fd597d5433058900630a350103b60b025a85a6850296050475d511a05684333a54015285a6600664e2744279a279027ae26a426ba26b61618280411106e497000000e780808f0000197186fca2f8a6f4caf0ceecd2e8d6e4dae0b2891306000232f80d46230cc10203b4090202e002e82af02ef461c003b589026307051083b409009305f5ff8e058d8113891500a10493058003330ab5026104854a17050000130b6589906001caa276027583b584ff946e829665ed08482ad803058401230ca1024c4803b509012eda033684ff0c6001ce631756019205aa95906563046601014621a08c618c61054632e02ee4033684fe833504ff01ce631756019205aa95906563046601014621a08c618c61054632e82eec0c6492052e95106508618a85029649e5c104130a8afc13048403e31b0af6b1a003ba890163080a0483b4090103b409001305faff12051181130915002104a104120a106001caa2760275833584ff946e829639e1906003b584ff8a8502960ded4104411ac104e31e0afc03b589006368a9002da0014903b589006371a90203b5090012092a99a27602758335090003368900946e829619c1054511a00145e6704674a6740679e669466aa66a066b09618280907588711c6e9765ffff9385d5a12d468287907588711c6e9765ffff938565a139468287411106e497f0ffffe78080740000411106e497f0ffffe780a0730000757106e5014730012948bd4821a89306f6ff13d547009a92a30f56fe0507368663fcf800aa879372f50013030003e3e002ff13037005e1bf13050008198d130610086370c5021765ffff930705a009462e85be8597000000e780e082aa60496182809305000897000000e78040660000757106e522e1a6fccaf8cef4d2f0d6ecdae8dee4e2e066fc6af86ef432892e8a014c814c814997f5000003bb25e897f5000083bb25e897f5000083b425e800690c612ef008652aec13058a002ae01765ffff130525972ae8294d22e40da03305b6000345f5ff5915133515002300a4006265146d02758296ee8c6311051213f5f90f631b051063758901e9a8636c890d33058941b3058a014146637fc50063022c0d81463386d50003460600630da6098506e319d5fe75a013867500937686ff3386b640ad8e93b6160013371600d98ea1c20146930605ff02676297b387c5009c6313c4f7ffa58fda9733747401e18f8defb307c7009c6313c4f7ffa58fda9733747401e18f95e34106e3f9c6fc31a83387d500034707006307a7038506e319d6fe930605ffe3f9c6fa6304c5062264b386c50083c606006386a6010506e319c5fe05a0b286e296138c1600e3f026f5d29603c50600e31ba5f38149e28de28a39a04a8c8549e68dca8a63872c030345040001c96265146d11460275c265829611ed33869a41b3059a01e39a9aed0145f1bd4a8c2264f9b7014511a00545aa600a64e6744679a679067ae66a466ba66b066ce27c427da27d49618280411106e41b8605009306000802c26376d6002302b100054671a01bd6b50019ee13d665001366060c2302c10093f5f50393850508a302b1000946ada01bd6050115e613d6c5001366060e2302c10013964503699213060608a302c10093f5f503938505082303b1000d462da81396b50275921306060f2302c1001396e502699213060608a302c100139645036992130606082303c10093f5f50393850508a303b10011464c0097000000e780e0d9a26041018280397106fc907594712ae032f836f4886d906994658c612af032ec36e82ee41765ffff930525810a85300097000000e78080b3e27021618280086117030000670063d5411106e408611b8605009306000802c26376d6002302b100054671a01bd6b50019ee13d665001366060c2302c10093f5f50393850508a302b1000946ada01bd6050115e613d6c5001366060e2302c10013964503699213060608a302c10093f5f503938505082303b1000d462da81396b50275921306060f2302c1001396e502699213060608a302c100139645036992130606082303c10093f5f50393850508a303b10011464c0097000000e78060caa26041018280397106fc90759471986d32f836f43af0906994658c61086132ec36e82ee42ae01755ffff930585710a85300097000000e780e0a3e27021618280357106ed22e926e54ae1cefcd2f8d6f42a840345050109c5833a04008544d5a0b2892e89033a840003654a03833a04009375450091e93336500163880a021755ffff9305e55e35a063960a0483358a0203350a02946d9755ffff9385855d094682961dc5814a854469a81755ffff9305655c83368a0203350a02946e05068296854441e103b689014a85d28502968da803254a038544a303910283350a0203368a022ee432e8930571022eec83250a0303068a0383360a0003378a0083370a0103388a01aaceaecc2300c10636f43af83efcc2e02800aae403b689011755ffff13052551aae82c104a85029619e9c6652665946d9755ffff9385655309468296aa8423089400850a233054012285ea604a64aa640a69e679467aa67a0d618280357106ed22e926e54ae1cefcd2f8d6f42a8403458500854a854419cd23049400a30454012285ea604a64aa640a69e679467aa67a0d6182803289ae89033a040003654a03834594001376450005e691cd83358a0203350a02946d9755ffff9385254b09468296854455f94e85d2850299aa846db785e183358a0203350a02946d9755ffff9385254905468544829659f503254a038544a303910283350a0203368a022ee432e8930571022eec83250a0303068a0383360a0003378a0083370a0103388a01aaceaecc2300c10636f43af83efcc2e02800aae41755ffff1305653faae82c104e85029915f9c6652665946d9755ffff9385a54109468296aa8439bf397106fc22f826f44af02a841c7508719c6f3a89b684829722e8230ca10002e4a30c01002800a6854a8697000000e78060db22658345810139c50544b9e5834591017d1513351500c264b335b0006d8d05c103c54403118901ed8c748870946d9755ffff9385153b05460544829611ed8c748870946d9755ffff9385a533054682962a8419a03334b0002285e2704274a274027921618280411106e497f0ffffe78020060000757106e5014730012948bd4831a89306f6ff9377f50f13d547009a92a30f56fe0507368663fbf8001373f50093020003e36f03fd93027003d9bf13050008198d130610086370c5021755ffff9307653209462e85be8597f0ffffe7804015aa60496182809305000897000000e780a0f80000757106e5014730012948bd4831a89306f6ff9377f50f13d547009a92a30f56fe0507368663fbf8001373f50093020003e36f03fd93027005d9bf13050008198d130610086370c5021755ffff9307452b09462e85be8597f0ffffe780200eaa60496182809305000897000000e78080f100001755ffff9306453809462e85b68517f3ffff6700232f397106fc22f826f42e848c752ae40870946d9755ffff938545384546829622ec2300a10202e8a30001021755ffff1306c53408082c0097000000e780a0c042658345010239c50544b9e5834511027d1513351500e264b335b0006d8d05c103c54403118901ed8c748870946d9755ffff9385552005460544829611ed8c748870946d9755ffff9385e518054682962a8419a03334b0002285e2704274a27421618280757106e5014730012948bd4821a89306f6ff13d547009a92a30f56fe0507368663fcf800aa879372f50013030003e3e002ff13037003e1bf13050008198d130610086370c5021755ffff9307c51809462e85be8597f0ffffe780a0fbaa60496182809305000897000000e78000df0000797106f422f026ec4ae84ee42a8404690865ae893309b640058d6363250308602695ce854a8697d00000e780a0f7ca9404e8a2700274e2644269a269456182802285a6854a8697000000e780c0000468f9b75d7186e4a2e026fc2e966368b6042a8408659314150063639600b284a14563e39500a14493c5f4fffd9119c5106032f0054632f42af811a002f428001410268697000000e780c003a265426581cdfd55fe158505630ab50009ed97b0ffffe7804002000008e004e4a6600664e2746161828097b0ffffe78020000000011106ec22e826e44ae03289aa8499cd2e84886605c18c6a91cd88624a8697b0ffffe780a0fc05e180e419a023b40400854521a8630409024a85a28597b0ffffe780c0f975d1814588e423b824018ce0e2604264a264026905618280228565f5e1b703e6450308619376060191ea1376060209ee0345050017f3ffff670063d10305050017030000670043d10305050017030000670063c903e6450308619376060189ea1376060219ea086117f3ffff670023ce086117f3ffff67008359086117030000670023e0411106e422e02a8411c96347040289c9228597b0ffffe78060f109a8054501a88545228597b0ffffe780c0ee19c9a285a26002644101828097b0ffffe78020f0000097b0ffffe780e0ee00005d7186e4a2e026fc4af84ef452f0ae898c750461006903b50902946d9755ffff9385a5f10546054982964ee42308a100a308010005c417050000930985f1138a140026ec28002c084e8697000000e78020a27d14d28465f40345010101ed22650c750871946d9755ffff938595f1054682962a894a85a6600664e2744279a279027a61618280797106f422f026ec4ae84ee42a8904690865058d2e84636fb50283390900894533859900636cb4007d148145228697d00000e780c0c3a2943385990023000500850423389900a2700274e2644269a269456182804a85a685228697000000e780e0008334090155bf5d7186e4a2e026fc2e966368b6042a8408659314150063639600b284a14563e39500a14493c5f4fffd9119c5106032f0054632f42af811a002f428001410268697000000e780c003a265426581cdfd55fe158505630ab50009ed97b0ffffe78060da000008e004e4a6600664e2746161828097b0ffffe78040d80000011106ec22e826e43284aa8499cd88660dc18c6a99cd8862228697b0ffffe78000d519ed85458ce431a823b40400854511a88545228597b0ffffe78040d27dd1814588e480e88ce0e2604264a26405618280411106e422e02a8408617d1508e005e90c70086c8c6182950870086511c5086c97b0ffffe78000cf087811c5087497b0ffffe78020ce08647d1508e409c5a2600264410182802285a2600264410117b3ffff670023cc5d7186e4a2e026fc4af84ef452f056ec83ba0501368a3289aa8963e3da00d28a806108687de1286c7d5610e8637c55010870106c98651c6d4e85b2854a86d286829761a08465306463edc400b386540163ee96082c683307b600636ec7086376d70208700c6c1074147c1c6d0a85268782970345010069e9a26563e8550f286c2ce824e426866367b50eb3b6c400918c33359500558d49e5338554016363950463e7a5080c7c63eca508b3059540639745090c74a6954a85528697d00000e78020af23b45901238009000868050508e8a6600664e2744279a279027ae26a616182801755ffff130565e611a81755ffff1305c5e529a01755ffff130525e5f14597f0ffffe780c00500001755ffff130575da9755ffff938665dbc1450a8689a01755ffff1305e5e89305f002d1bf1755ffff1305f5ea93052003d9b7528597000000e780408b00001755ffff1305e5059755ffff938605dd9305b0021306710197f0ffffe780c01a00001755ffff1305a5df71b71755ffff1305c5e09305e00241b7034505000e051756ffff130606392a969756ffff9386663d369598751062146188711c6fb6858287411110650c69b29563edc50008611069fd568582637dd60028616369b502410182801755ffff1305c5aea14535a01755ffff130505d19755ffff938605d2e145300097f0ffffe780001200001755ffff130595e19305600297f0ffffe780a0f50000797106f422f0aa8502c2280050009146114497000000e78020de0345810011e942656319850203654100a2700274456182801755ffff130585f69755ffff9386a5cd9305b0021306f10197f0ffffe780600b00001755ffff130555ddb54597f0ffffe78020ef0000411106e497000000e78040f98d4563f7a50009817d15a260410182801755ffff130525dbb94597f0ffffe78020ec0000197186fca2f8a6f4caf0ceecd2e8d6e4dae05efc03bb050003370b00806594692a89130517002330ab0065c95ae409072330eb007dc3b28a36f85af02e8597000000e780a0f29305440063ea850caa892ef4081097000000e780c0f763ffaa02aa84938b1a0013952b002295636e850a2af4081097000000e78040ef2a8a63999b02330544016366850a2ae863f649051755ffff130565dfc1a015452304a900233009005a8597000000e78000c6b1a08a0a33858a002105636285082af4081097000000e78080eab305440163ed8506aa892ee8636e4507338549412aec280097000000e78060e26265c26522662338a9002334b9002330c9005a8597000000e780a0c0e6704674a6740679e669466aa66a066be27b09618280000000001755ffff130585d60da81755ffff1305e5d525a01755ffff130545d539a81755ffff1305a5d411a81755ffff130505d429a01755ffff130565d39305b00297f0ffffe780c0d50000797106f422f0906118629465050718e20dcf2a841385460032e4636ad5022ae82e8597000000e78000de2aec280097000000e78020d76265c265226608e80ce410e0a270027445618280000000001755ffff130525cd9305b00297f0ffffe78080cf0000397106fc22f826f42a8402e408083000a146a144a28597000000e780c0b70345010105e16265631f9502a264086097000000e780e0b02685e2704274a274216182801755ffff130565cf9755ffff938685a69305b0021306710297f0ffffe78040e400001755ffff1305e5b7b94597f0ffffe78000c80000397106fc22f826f42a84a307010008081306f10085468544a28597000000e78000b0034501010de16265631095048304f100086097000000e78000a92685e2704274a274216182801755ffff130585c79755ffff9386a59e9305b0021306710297f0ffffe78060dc00001755ffff1305c5b1b54597f0ffffe78020c000005d7186e4a2e026fc4af8ae842a898c69054632e002e402e889c90a8597000000e780408f0266426411a001442808a685a28697000000e780a0a6034581011de5027563168504c2652266826688602338b9002334c9002330d900a6600664e27442796161170300006700239e1755ffff130565bd9755ffff938685949305b0021306f10297f0ffffe78040d200001755ffff130575a8c94597f0ffffe78000b60000011106ec22e826e49c692a84637df700b384e74063e3d400b684b306970063ede60263f7d7001545a300a400054531a8998e639dd4028c61ba953285268697c00000e7808056014504e42300a400e2604264a264056182801755ffff1305a58ef14597f0ffffe78040af00002685b68597f0ffffe780c03700005d7186e4a2e026fc4af84ef452f02e8483b905012a896145a14597a0ffffe780806159c1aa84086888e8086488e4086088e0054a52e402e802ec1314ba002800a28597f0ffffe780207b13050006a14597a0ffffe780205e21c923304501233445012338050004ed9755ffff9385859a0cf1a2650cf5c2650cf9e2650cfd23303505233405042338050420ed23340900233839012330a900a6600664e2744279a279027a6161828097a0ffffe780a05a00000c6591c5086117a3ffff670023588280397106fc22f826f44af09376f60f1307f00f2a89638fe6041b04160002ec02e802e402e0131584036d9113060002098e8a84aa94aa95268597c00000e78020431375740009c9838504007d563315a6006d8d2380a4008a85130600024a8597c00000e780c040e2704274a274027921618280130600024a858145e2704274a2740279216117c30000670083312a860345050283c605023337d500358d3335a000b306e040558d0de5fd057d06815695c20345060003c70500b337e500398d3335a0003307f040598dfd157d16850665d18280014582805d7186e4a2e026fc4af8ae84806590612a892800a28597e0ffffe780c0020345810019c5426529e109452300a90029a805040dc09305910080e4130610024a8597c00000e7804035a6600664e2744279616182801755ffff1305c58ef14597f0ffffe780608e000097e0ffffe780801d0000306115ce14610c653337d00093b715007d8f7d1630e115c7106d0c699306050109c683b505227d166dfe0146014723b4060023b00600854614e10ce531a08145b1a8b5ca1869106d83d6a5216374d600ae8621a883b60521a1c603d6852183d7a6210507b685e377f6fe1308160001cf0e083698833708227d1701c783b70722e5bf014811a0b68793050003b305b602b6951ce523380500233c05012e8582801755ffff130505809305b00297f0ffffe780608200001745ffff1305a57eedb7411106e413050022c14597a0ffffe780e03501c5a2604101828097a0ffffe780e0360000411106e413050028c14597a0ffffe780a03301c5a2604101828097a0ffffe780a03400001d7186eca2e8a6e4cae04efc52f856f45af05eec62e866e46ae03e893a8ab689b28aae8b2a84035ca52193841500139b55002a9b139d4500b30cbc40637b9c00130600025a85d68597c00000e780201d81a013955400229513965c00da8597c00000e780a060130600025a85d68597c00000e780c01a13050416b305a50113964400329513964c0097c00000e780005e930a1c00229d23344d1723303d1793092c00130a042213852b00139b3400637c3501b3056a010e05529513963c0097c00000e780a05a5a9a23302a01231d542163f434038e0ba29b13858b22b305804109461461239c9620850423b88620b38695002105e397c6fee6604664a6640669e279427aa27a027be26b426ca26c026d256182800358a5212e86814593125800aa929303f5011303f601054e63055504938815001305050201579a869e8715cf83ce060003c6070033bfce0033c6ce00b33ec0003306e0413366d601fd17fd16050771de1376f60f631ac60193830302c685e31f55fac28511a0014e72858280457186e7a2e326ff4afb4ef752f356ef5aeb5ee762e3e6feeafaeef62e8a83bb050083b90501b28a2a8b03d9ab21139559005e9583459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18d2ef483451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2ef083459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2eec83451500034605008346250003473500a205d18dc2066207d98ed58d034655008346450003476500834775002206558e4207e2075d8f598e0216d18d2ee8938c190093955c00de9513c6f9ff330426011316540097c00000e780603a93850b16139549002e950465033c050013964c00b2951316440097c00000e78040387d3913150903239d2b21033a8a0041919545637bb51a2819de85528697000000e780601f6a7556e026e405cd85456317b5068001080113068003a28597c00000e78020ef6a65aa750355a52183d5a5212e950505b1456376b50408180c01014605a88001a80013068003a28597c00000e78020ec0675c6750355a52183d5a5212e950505b1456372b5040818ac000546ce8697000000e780e04e99a80e65ae650da0081a13068003a28597c00000e78040e8081a854597000000e780401c3665d6652af82efccee025a0081a13068003a28597c00000e780c0e5081a854597000000e780a078766596752af82efce6e0c27b627a03b60b21866971c613041a00930a010c914c314d954d05498354a62163eb9c0a2819b285228697000000e780800f6a751dcd631b2509a81913068003d68597c00000e780c0df526592750355a52183d5a5212e950505636ea503b3859d40a81997000000e780601201465df69da0a81913068003d68597c00000e78040dc526592750355a52183d5a5212e9505056373a503081a13068003d68597c00000e78000da081a97100000e780009a2a862e8425f605a0b3859d40a81997000000e780a06b014631fa31a089e4054582652380a500a264227582756266c266233cab002338bb002334cb002330db0023308b0323349b0223387b03233c4b0323303b05be601e64fa745a79ba791a7afa6a5a6bba6b1a6cf67c567db67d7961828083b605219dc683d78521130816009dc71387f7ff93173700b69783b707222330050014e52338050118ed1cf110f50cf92da00ce510e989450ce1828003d7a62119cf03b7862285471ce114e523380501233c05000cf110f518f910fd828097e0ffffe780a0b60000317106fd22f926f54af14eed52e956e55ae1defce2f8e6f4eaf0eeec6383052a2e892a8a833b850183d5ab21338425012d45636e85282ef4033b8a020355ab21636e252933052541239d8b202ae4231dab20930af9ff93945a0093090b1613954a002ae84e9583350a01833d0a00106532f008612aec139555006e959205ae9d83459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18daee483451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18daee083459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2efc83451500034605008346250003473500a205d18dc206620703465500d98ecd8e83454500220603476500834775004d8e268cb3059b004207e2075d8f598e0216558e32f81306000297c00000e78000f803bd0d1683bc8d16626523b0ad16027523b4ad16a28da274139554005e950c181306000297c00000e78060b013840b16139544002295233495018504b3859d402330a501639cba10139554005e95da85628697c00000e78080ad139544002295ce85426697c00000e78060ac93155900da95226c13165c005a8597c00000e780e0ef93154900ce9513164c004e8597c00000e780a0ee83350a0203350a03adcd79c113040b22139534005e951305052293193900a2854e8697c00000e78020a7b305340113163c002106228597c00000e780c0eaa27c63f0bc038e0cde9c13858c220c61239c9520850423b875217d192105e31809fe7d556301ac020145050c0c601306150023b86521239ca52021043285e317ccfe11a039e5ea704a74aa740a79ea694a6aaa6a0a6be67b467ca67c067de66d296182801745ffff1305c512ed4505a81745ffff1305d51b930520030da01745ffff1305151e11a81745ffff1305b50a29a01745ffff130535179305800297e0ffffe78080f60000317106fd22f926f54af14eed52e956e55ae1defce2f8e6f4eaf0eeec806d035da4216a8701c698750357a721636cd72832f036f42af883ba850203dcaa21930b1d0033868b012d456365c528846188652ae803b9050188712aec03dba42132e4231dc42013155900269583459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18daee883451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18daee483459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18daee083451500034605008346250003473500a205d18dc2066207d98ed58d034655008346450003476500834775002206558e4207e2075d8f598e0216d18d2efc930d190093955d00a6959349f9ffda991396590097c00000e78060c813155d0022952c181306000297c00000e780408213955b00229513165c00d68597c00000e780008193850416131549002e95033a0500833c850013964d00b2951396490097c00000e780a0c31305041693154d00aa9523b4950123b0450193850a1613964b00329513164c0097b00000e780407c9385042213953d002e950e09ca95c1051396390097c00000e78060bf63f06d032699130589220c6113861d0023b89520239cb5212105b28de317cbfe0395a4217d358545239da420426563f3a50413953b0022951305052293850a2213163c00210697b00000e780a07522656372ad02050c0e0d229d13058d22de851061231cb6208505233886207d1c2105e3180cfe027593341500568597a0ffffe7802083fd1433f57401a2752e95c27580e1626690e588e9ea704a74aa740a79ea694a6aaa6a0a6be67b467ca67c067de66d296182801745ffff1305b5f19305100939a01745ffff1305e5f99305a00297e0ffffe78000c80000717106f522f126ed4ae94ee552e1d6fcdaf8def4e2f0e6eceae8eee4638605262e8b2a890075835ca421e6952d456363b526033c89018354ac2163e46427338d6441231dac212ee4231db42013155b00229513965c00a28597c00000e780c0ab9309041613154b004e9513964c00ce8597c00000e78040aa930b1d00b38a74411305fbff6396aa2293955b00e295139a5a002285528697b00000e780006393040c1693954b00a695920a4e85568697b00000e780806113154d00269583350901833d0900106532ec08612ae8139555006e959205ae9d83459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18d2efc83451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2ef883459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2ef483451500034605008346250003473500a205d18dc20662070346550083474500d98ecd8e22065d8e034765008347750093155d00e2954207e2075d8f598e0216558e32f01306000297c00000e780c09303bd0d1683b48d16426523b0ad16626523b4ad16330544010c101306000297b00000e780804cd69923b4990023b0a9018335090203350903a1c945c1930404220e0b3385640113963c002106a68597c00000e780608e8e0be29b93850b2226855a8697b00000e780404881452265050590609386150023388620231cb620a104b685e317d5fe11a029e9aa700a74ea644a69aa690a6ae67a467ba67b067ce66c466da66d4d6182801745ffff130585b7ed4515a81745ffff130575b8930530031da01745ffff1305c5ba9305700221a81745ffff130535af29a01745ffff1305b5bb9305800297e0ffffe780009b0000357106ed22e926e54ae1cefcd2f8d6f4daf0deece2e8e6e4eae06efc033a850183398502835aaa2103dba92113841a0033066401ad4563e1c526033d0500833c050108652ae8035cad2132e4231dca2013955c006a9583459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18d2ef883451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2ef483459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2ef083451500034605008346250003473500a205d18dc2066207d98ed58d034655008346450003476500834775002206558e4207e2075d8f598e0216d18d2eec93841c0093955400ea9593cdfcffe29d13965d0097b00000e780206e13955a0052952c081306000297b00000e780002813155400529513165b00ce8597b00000e780c02693050d1613954c002e9503390500833b850013964400b29513964d0097b00000e780606913050a1693954a00aa9523b4750123b025019385091613164400329513164b0097b00000e780002293050d22139534002e958e0ce695c10513963d0097b00000e780206563f08403ea9c13858c220c611386140023b8a521239c95202105b284e317ccfe0315ad217d358545231dad20c26463f29504131534005295130505229385092213163b00210697b00000e780601b226563f1aa02050b8e0ad29a13858a220c61239c8520050423b845217d1b2105e3180bfe4e859790ffffe78060296a85a685ea604a64aa640a69e679467aa67a067be66b466ca66c066de27d0d6182801745ffff130505a29305a00297d0ffffe78020700000411106e413058072a1459790ffffe780402401c5a260410182809790ffffe78040250000411106e413058078a1459790ffffe780002201c5a260410182809790ffffe780002300001d7186eca2e8a6e4cae04efc52f856f45af05eec62e866e43a89b689328a2e8b2a84835b655b1305855b938415009605da95b30ab500338c6b4163fb9b00130610025685d28597b00000e780a00ba9a09395540026952e9513165c006296d68597b00000e780e04e130610025685d28597b00000e78000091305840013064008b305cb02aa95b386c40236953306cc0297b00000e780e04b138a1b00130540083305ab022295210513064008ce8597b00000e780200593892b00930a847213052b00939c3400637c3501b3859a010e05569513163c0097b00000e7808047e69a23b02a01231b445b63f334030e0b229b13050b73b305704109461461239a965a850480e2b38695002105e398c6fee6604664a6640669e279427aa27a027be26b426ca26c25618280397106fc22f826f44af04eec52e856e48359655b2e8a9305855b93945900ce947d54054995c4938a1502528597f0ffffe780e0bc9384f4fd1375f50f0504d685e30225ff9305f00f6305b500014911a04e844a85a285e2704274a2740279e269426aa26a21618280130101ce233c1130233881302334913023302131233c312f2338412f2334512f2330612f233c712d2338812d2334912d2330a12d233cb12b2e8c83bb050003bb05013289aa8903da6b5b13848b5b13155b005a95b30ca400a80b13061002e68597b00000e78000f1930a1b0093955a005694a2951345fbffb3044501139654002696668597b00000e780a033930c400833059b033384ab00130d84001305911f13064008ea8597b00000e780a0ec9305c408338694036a8597b00000e78060301b05faff239bab5a033a8c004215135405032811ac0b1306500a97b00000e78060e90a852c111306500a97b00000e78060e81545637da41a2811de85528697000000e78060202a7505cd85456317b5060019081313068003a28597b00000e78060e57a75be650355655b83d5655b2e950505b1456376b504880a0c13014605a80019a81213068003a28597b00000e78060e21a65da650355655b83d5655b2e950505b1456372b504880aac120546da8697000000e780004ca9a84a75ea750da0a80b13068003a28597b00000e78080dea80b854597000000e780601d5e75fe75aaeaaeeedaf235a0a80b13068003a28597b00000e78000dca80b854597000000e780a06b0335012083358120aaeaaeeed6f2d66b766a03b60b00167b69ca93041a00930a010b914d314c954c054d0354665b63ee8d0a2811b285268697000000e78080102a7529c1631fa509080513068003d68597b00000e780c0d5033581298335812a0355655b83d5655b2e95050563608505b3858c40080597000000e780001301464df6a5a0080513068003d68597b00000e78000d2033581298335812a0355655b83d5655b2e95050563738503a80b13068003d68597b00000e78080cfa80b97100000e78020882a86ae8425f239a8b3858c40080597000000e780e05d014631f629a001e405452300a9008a851306500a4e8597b00000e780a0cb23b4790b23b8490b23bc690b833081310334013183348130033901308339812f033a012f833a812e033b012e833b812d033c012d833c812c033d012c833d812b13010132828094619dc683d7455b130816009dc71387f7ff93173700b69783b787722330050014e52338050118ed1cf110f50cf92da00ce510e989450ce1828003d7665b19cf03b7067385471ce114e523380501233c05000cf110f518f910fd828097d0ffffe780c0ab0000130101d92334112623308126233c9124233821252334312523304125233c5123233861232334712323308123233c91212338a1212334b121638505242e89aa8b033d850103546d5bb304b4002d456360952422ec83bc8b0203d56c5b63602525330a2541231b9d5a239b4c5b930df9ff93898c5b13955d006e952ae4338ba900938a8c0013044008b3858d022ee8d69528101306400897b00000e78000b703b50b0183b50b0013165500b386a500369626f09304865b330585022e95130c8500081913061002a68597b00000e780e0b3130610022685da8597b00000e780c0f79304110d130640082685e28597b00000e780a0b12c1013064008628597b00000e780a0b0a80a0c191306100297b00000e780a0af080313064008a68597b00000e780a0ae130b8d5b626c13155c00b3058b012e95ac0a1306100297b00000e780c0ac93048d0033058c0226950c031306400897b00000e78040ab13041c000275018d6392ad1413155400229b5a95ce85226697b00000e78040a9130b4008330564032695d685426697b00000e780e0a7131559004a95b385a90013165a0052964e8597b00000e78020ebb3056903d69533066a03568597b00000e780e0e983b50b0203b50b03c1c165c5d28a93848c72131534006a951305857293193900a6854e8697b00000e78040a2b385340113163a002106268597b00000e780e0e502756371ac02131a3c006a9a13050a730c61239a855a050423b0a5017d192105e31809fe7d556382aa02814513851a0090609386150023309601231ab65aa104b685e317d5fe11a02de58330812603340126833481250339012583398124033a0124833a8123033b0123833b8122033c0122833c8121033d0121833d81201301012782801735ffff1305e50bed4505a81735ffff1305f514930520030da01735ffff1305351711a81735ffff1305d50329a01735ffff130555109305800297d0ffffe780a0ef0000697106f622f226ee4aea4ee652e2d6fddaf9def5e2f1e6edeae9eee583bd850103dc6d5b628701c698750357675b636ad71e32f036f42af883ba850283dc6a5b130b1c0033069b012d456363c51e846188652ae888712aec83b9050183db645b32e4239bcd5a1384845b139559004e95330da400880013061002ea8597b00000e780408c13891900931559004a94a29513caf9ff5e9a52fc13165a0052966a8597b00000e780e0ce13848d5b13155c00b30584012e958c001306100297b00000e780408893858a5b13155b005a94229513965c00669697b00000e780a086130d40083385a9033384a400628a5a8c668bd68c930a8400880013064008d68597b00000e78020849305c40862753306a5035685e68ada8c628b97b00000e78060c713848d003305aa0322958c001306400897b00000e780008193858a003305ac0322953386ac0397a00000e780a07f93858472131539002e958e09ce95c10562760e0697b00000e780c0c2637f7901a699138509730c611306190084e1239a255b21053289e398cbfe0395645b7d358545239ba45a426563f4a50413153b006e951305857293858a7213963c00210697a00000e780207922656373aa02850c131c3a006e9c13050c73da851061231ab65a85052330b601fd1c2105e3980cfe02751334150056859790ffffe78080867d1433756401a2752e95c27523b0b501626690e588e9b2701274f2645269b269126aee7a4e7bae7b0e7cee6c4e6dae6d556182801735ffff1305f5f49305100939a01735ffff130525fd9305a00297d0ffffe78040cb0000130101d92334112623308126233c9124233821252334312523304125233c5123233861232334712323308123233c91212338a1212334b121638705202e8caa8b0075035d645bea952d456364b52003bb8b01835a6b5b63e58a21338a8a41231b4b5b2ee8231bb45a1309845b13155c0062954a9513165d006a96ca8597b00000e780c0ac93098400930c400833059c034e9533069d03ce8597b00000e78000ab930d1a00b384ba411305fcff6391a41cda8a130b8b5b93955d003305bb01aa95139554003306950032f04a8597a00000e780e06256e4a10ab3859d03d6953386940332ec4e8597a00000e780406113155a00529b2a9bb3059a03d69528101306400897a00000e780805f03b50b0183b50b0013165500b386a50036969304865b330595032e95930c8500081913061002a68597a00000e780805c130610022685da8597b00000e78060a09304110d130640082685e68597a00000e780405a2c1013064008668597a00000e7804059a80a0c191306100297a00000e7804058080313064008a68597a00000e780405702754a95ac0a1306100297a00000e780205662654e950c031306400897a00000e780005583b50b0203b50b03a1c955cd930484720e0c3385840113163d002106a68597b00000e78080978e0d2265aa9d93858d722685628697a00000e780405181454265050590609386150000e2231ab65aa104b685e318d5fe11a03de58330812603340126833481250339012583398124033a0124833a8123033b0123833b8122033c0122833c8121033d0121833d81201301012782801735ffff1305e5beed4515a81735ffff1305d5bf930530031da01735ffff130525c29305700221a81735ffff130595b629a01735ffff130515c39305800297d0ffffe78060a200006d7106e622e2a6fdcaf9cef5d2f1d6eddae9dee5e2e166fd6af96ef5033a850183398502035b6a5b83db695b13041b0033067401ad4563ebc51a833c05000c652eec833d050103dd6c5b32e0231bca5a13898c5b13955d006e95b30aa900081013061002d68597a00000e780604093841d00939554002699ca9513c9fdff6a99131659004a96568597b00000e7802083930a8a5b13155b00b3856a012e950c101306100297a00000e780803c9385895b13155400a29a569513965b005e9697a00000e780e03a130c400833858d03b38aac005ee4ce8b93898a00081013064008ce8597a00000e780a0389385ca08330689034e8597a00000e780607c93098a005ae833058b034e950c101306400897a00000e780e035de8a93858b00a26b330584034e9533868b0397a00000e780403493858c72139534002e958e0dee95c1051316390097a00000e780607763f0a403e69d13850d730c611386140023b09501239a955a2105b284e317cdfe03956c5b7d358545239bac5ae264426b63f295041315340052951305857293858a7213963b00210697a00000e780802d02656371ab02850b0e0b529b13050b730c61239a855a050423b04501fd1b2105e3980bfe56859780ffffe780803b6685a685b2601264ee744e79ae790e7aee6a4e6bae6b0e6cea7c4a7daa7d516182801735ffff130525b49305a00297d0ffffe78040820000130101dc233c1122233881222334912223302123233c3121233841212334512123306121deffe2fbe6f7eaf3eeefd54bae8a63f575052a8c094563e9aa0005466285d68597300000e78040e98330812303340123833481220339012283398121033a0121833a8120033b0120fe7b5e7cbe7c1e7dfe6d130101248280b68cb2892afc930d7113054d0545aae856f8627c1b850c0019e16f20f00613751d0019e16f10b07d466813db2a0013171b00b308670113051003637955231303fbff93021b0013166b00629603459601834586018346a6018347b60122054d8dc206e207dd8e558d8345d6018346c6018347e6018344f601a205d58dc207e204c58fdd8d82154d8d2af90345160183450601834626018347360122054d8dc206e207dd8e558d83455601834646018347660183447601a205d58dc207e204c58fdd8d82154d8d2af503459600834586008346a6008347b60022054d8dc206e2078345d6008344c600dd8e558da205cd8c8346e6008347f60093156300e295c206e207dd8ec58e8216558d2af1034516008346060083472600834436002205558dc207e204c58f5d8d83465600834746008344660003467600a206dd8ec2046206458e558e0216518d2aed03c5950103c6850183c6a50183c7b5012205518dc206e207dd8e558d03c6d50183c6c50183c7e50183c4f5012206558ec207e204c58f5d8e0216518d2afa03c5150103c6050183c6250183c735012205518dc206e207dd8e558d03c6550183c6450183c7650183c475012206558ec207e204c58f5d8e0216518d2af603c5950003c6850083c6a50083c7b5002205518dc206e207dd8e558d03c6d50083c6c50083c7e50083c4f5002206558ec207e204c58f5d8e0216518d2af203c5150003c6050083c6250083c735002205518dc206e207dd8e558d03c6550083c6450083c7650083c575002206558ec207e205dd8dd18d82154d8d2aee01559305710b6e8605c583c60500834706007d16fd150505e388f6feb3b3f60063f9f6009a875a8331a081436f10c0168143da8713956200629503469501834685018344a5010344b5012206558ec2046204458c418e8346d5018344c5010344e5018345f501a206c58e4204e205c18dd58d8215d18d2ef983451501034605018346250183443501a205d18dc206e204c58ed58d034655018346450183446501034475012206558ec2046204458c418e0216d18d2ef583459500034685008346a5008344b500a205d18dc206e2040346d5000344c500c58ed58d2206518c8346e5008344f500139667006296c206e204c58ec18e8216d58d2ef183451500834605008344250003443500a205d58dc2046204458cc18d83465500834445000344650003457500a206c58e42046205418d558d02154d8d2aed03459601834586018346a6018344b60122054d8dc206e204c58e558d8345d6018346c6018344e6010344f601a205d58dc2046204458cc18d82154d8d2afa0345160183450601834626018344360122054d8dc206e204c58e558d83455601834646018344660103447601a205d58dc2046204458cc18d82154d8d2af603459600834586008346a6008344b60022054d8dc206e204c58e558d8345d6008346c6008344e6000344f600a205d58dc2046204458cc18d82154d8d2af20345160083450600834626008344360022054d8dc206e204c58e558d83455600834646008344660003467600a205d58dc2046206458ed18d82154d8d2aee01551306710b130471130dc183440600834604007d147d160505e388d4fe63e3d400be8233b5d400aa93968713956700629583459501034685018346a5018344b501a205d18dc206e204c58ed58d0346d5018346c5018344e5010344f5012206558ec2046204458c418e0216d18d2ef983451501034605018346250183443501a205d18dc206e204c58ed58d034655018346450183446501034475012206558ec2046204458c418e0216d18d2ef583459500034685008346a5008344b500a205d18dc206e2040346d5000344c500c58ed58d2206518c8346e5008344f500131663006296c206e204c58ec18e8216d58d2ef183451500834605008344250003443500a205d58dc2046204458cc18d83465500834445000344650003457500a206c58e42046205418d558d02154d8d2aed03459601834586018346a6018344b60122054d8dc206e204c58e558d8345d6018346c6018344e6010344f601a205d58dc2046204458cc18d82154d8d2afa0345160183450601834626018344360122054d8dc206e204c58e558d83455601834646018344660103447601a205d58dc2046204458cc18d82154d8d2af603459600834586008346a6008344b60022054d8dc206e204c58e558d8345d6008346c6008344e6000344f600a205d58dc2046204458cc18d82154d8d2af20345160083450600834626008344360022054d8dc206e204c58e558d83455600834646008344660003467600a205d58dc2046206458ed18d82154d8d2aee01551306710b9304711315c10344060083c60400fd147d160505e308d4fe6363d4003e833335d400aa931a8b11a03e8b9304f7ff9362170013156700629583459501034685018346a5018347b501a205d18dc206e207dd8ed58d0346d5018346c5018347e5010344f5012206558ec2076204c18f5d8e0216d18d2ef983451501034605018346250183473501a205d18dc206e207dd8ed58d034655018346450183476501034475012206558ec2076204c18f5d8e0216d18d2ef583459500034685008346a5008347b500a205d18dc206e2070346d5000344c500dd8ed58d2206518c8346e5008347f500139664006296c206e207dd8ec18e8216d58d2ef183451500834605008347250003443500a205d58dc2076204c18fdd8d83465500834745000344650003457500a206dd8e42046205418d558d02154d8d2aed03459601834586018346a6018347b60122054d8dc206e207dd8e558d8345d6018346c6018347e6010344f601a205d58dc2076204c18fdd8d82154d8d2afa0345160183450601834626018347360122054d8dc206e207dd8e558d83455601834646018347660103447601a205d58dc2076204c18fdd8d82154d8d2af603459600834586008346a6008347b60022054d8dc206e207dd8e558d8345d6008346c6008347e6000344f600a205d58dc2076204c18fdd8d82154d8d2af20345160083450600834626008347360022054d8dc206e207dd8e558d83455600834646008347660003467600a205d58dc20762065d8ed18d82154d8d2aee01551306710b9306711315c18347060003c40600fd167d160505e38887fe33b58700aa9363f58700a686ba8411a0ba8613956200629583459501034685010347a5018347b501a205d18d4207e2075d8fd98d0346d5010347c5018347e5010344f5012206598ec2076204c18f5d8e0216d18d2ef983451501034605010347250183473501a205d18d4207e2075d8fd98d034655010347450183476501034475012206598ec2076204c18f5d8e0216d18d2ef583459500034685000347a5008347b500a205d18d4207e2070346d5000344c5005d8fd98d2206518c0347e5008347f5001396660062964207e2075d8f418f0217d98d2ef183451500034705008347250003443500a205d98dc2076204c18fdd8d0347550083474500034465000345750022075d8f42046205418d598d02154d8d2aed03459601834586010347a6018347b60122054d8d4207e2075d8f598d8345d6010347c6018347e6010344f601a205d98dc2076204c18fdd8d82154d8d2afa0345160183450601034726018347360122054d8d4207e2075d8f598d83455601034746018347660103447601a205d98dc2076204c18fdd8d82154d8d2af603459600834586000347a6008347b60022054d8d4207e2075d8f598d8345d6000347c6008347e6000344f600a205d98dc2076204c18fdd8d82154d8d2af20345160083450600034726008347360022054d8d4207e2075d8f598d83455600034746008347660003467600a205d98dc20762065d8ed18d82154d8d2aee01551306710b130771130dc103440600834707007d177d160505e308f4fe6363f400b6823335f400aa93968613956600629583459501034685010347a5018347b501a205d18d4207e2075d8fd98d0346d5010347c5018347e5010344f5012206598ec2076204c18f5d8e0216d18d2ef983451501034605010347250183473501a205d18d4207e2075d8fd98d034655010347450183476501034475012206598ec2076204c18f5d8e0216d18d2ef583459500034685000347a5008347b500a205d18d4207e2070346d5000344c5005d8fd98d2206518c0347e5008347f5001396640062964207e2075d8f418f0217d98d2ef183451500034705008347250003443500a205d98dc2076204c18fdd8d0347550083474500034465000345750022075d8f42046205418d598d02154d8d2aed03459601834586010347a6018347b60122054d8d4207e2075d8f598d8345d6010347c6018347e6010344f601a205d98dc2076204c18fdd8d82154d8d2afa0345160183450601034726018347360122054d8d4207e2075d8f598d83455601034746018347660103447601a205d98dc2076204c18fdd8d82154d8d2af603459600834586000347a6008347b60022054d8d4207e2075d8f598d8345d6000347c6008347e6000344f600a205d98dc2076204c18fdd8d82154d8d2af20345160083450600034726008347360022054d8d4207e2075d8f598d83455600034746008347660003467600a205d98dc20762065d8ed18d82154d8d2aee01551306710b1307711315c183470600034407007d177d160505e38887fe63e38700b68433b58700aa93268711a036871383f8ff9382180013956800629583459501034685018346a5018347b501a205d18dc206e207dd8ed58d0346d5018346c5018347e5018344f5012206558ec207e204c58f5d8e0216d18d2ef983451501034605018346250183473501a205d18dc206e207dd8ed58d034655018346450183476501834475012206558ec207e204c58f5d8e0216d18d2ef583459500034685008346a5008347b500a205d18dc206e2070346d5008344c500dd8ed58d2206d18c8346e5008347f500131663006296c206e207dd8ec58e8216d58d2ef183451500834605008347250083443500a205d58dc207e204c58fdd8d83465500834745008344650003457500a206dd8ec2046205458d558d02154d8d2aed03459601834586018346a6018347b60122054d8dc206e207dd8e558d8345d6018346c6018347e6018344f601a205d58dc207e204c58fdd8d82154d8d2afa0345160183450601834626018347360122054d8dc206e207dd8e558d83455601834646018347660183447601a205d58dc207e204c58fdd8d82154d8d2af603459600834586008346a6008347b60022054d8dc206e207dd8e558d8345d6008346c6008347e6008344f600a205d58dc207e204c58fdd8d82154d8d2af20345160083450600834626008347360022054d8dc206e207dd8e558d83455600834646008347660003467600a205d58dc20762065d8ed18d82154d8d2aee01551306710b9304711315c18346060083c70400fd147d160505e388f6fe33b5f600aa9363f5f6001a86468311a0468613956200629583459501834685018347a5018344b501a205d58dc207e204c58fdd8d8346d5018347c5018344e5010344f501a206dd8ec2046204458cc18e8216d58d2ef983451501834605018347250183443501a205d58dc207e204c58fdd8d83465501834745018344650103447501a206dd8ec2046204458cc18e8216d58d2ef583459500834685008347a5008344b500a205d58dc207e2048346d5000344c500c58fdd8da206c18e8347e5000344f50093146600e294c2076204c18fdd8e8216d58d2ef183451500834605008347250003443500a205d58dc2076204c18fdd8d83465500834745000344650003457500a206dd8e42046205418d558d02154d8d2aed03c5940183c5840183c6a40183c7b40122054d8dc206e207dd8e558d83c5d40183c6c40183c7e40103c4f401a205d58dc2076204c18fdd8d82154d8d2afa03c5140183c5040183c6240183c7340122054d8dc206e207dd8e558d83c5540183c6440183c7640103c47401a205d58dc2076204c18fdd8d82154d8d2af603c5940083c5840083c6a40083c7b40022054d8dc206e207dd8e558d83c5d40083c6c40083c7e40003c4f400a205d58dc2076204c18fdd8d82154d8d2af203c5140083c5040083c6240083c7340022054d8dc206e207dd8e558d83c5540083c6440083c7640083c47400a205d58dc207e204c58fdd8d82154d8d2aee01559304710b130471130dc183c70400834604007d14fd140505e388d7fe63e3d700b28233b5d700aa93168613156600629583459501834685018347a5018344b501a205d58dc207e204c58fdd8d8346d5018347c5018344e5010344f501a206dd8ec2046204458cc18e8216d58d2ef983451501834605018347250183443501a205d58dc207e204c58fdd8d83465501834745018344650103447501a206dd8ec2046204458cc18e8216d58d2ef583459500834685008347a5008344b500a205d58dc207e2048346d5000344c500c58fdd8da206c18e8344e5000344f50093176300e297c2046204458cc18e8216d58d2ef183451500834605008344250003443500a205d58dc2046204458cc18d83465500834445000344650003457500a206c58e42046205418d558d02154d8d2aed03c5970183c5870183c6a70183c4b70122054d8dc206e204c58e558d83c5d70183c6c70183c4e70103c4f701a205d58dc2046204458cc18d82154d8d2afa03c5170183c5070183c6270183c4370122054d8dc206e204c58e558d83c5570183c6470183c4670103c47701a205d58dc2046204458cc18d82154d8d2af603c5970083c5870083c6a70083c4b70022054d8dc206e204c58e558d83c5d70083c6c70083c4e70003c4f700a205d58dc2046204458cc18d82154d8d2af203c5170083c5070083c6270083c4370022054d8dc206e204c58e558d83c5570083c6470083c4670083c77700a205d58dc204e207c58fdd8d82154d8d2aee01559307710b9304711315c103c4070083c60400fd14fd170505e308d4fe6363d40032833335d400aa939a8811a0b28813156700629503469501834685018347a5018344b5012206558ec207e204c58f5d8e8346d5018347c5018344e5010344f501a206dd8ec2046204458cc18e8216558e32f9034615018346050183472501834435012206558ec207e204c58f5d8e83465501834745018344650103447501a206dd8ec2046204458cc18e8216558e32f503469500834685008347a5008344b5002206558ec207e2048346d5000344c500c58fd18fa206c18e8344e5000344f50013166b006296c2046204458cc18e8216dd8e36f183461500834705008344250003443500a206dd8ec2046204458cc18e83475500834445000344650003457500a207c58f42046205418d5d8d0215558d2aed03459601834686018347a6018344b6012205558dc207e204c58f5d8d8346d6018347c6018344e6010344f601a206dd8ec2046204458cc18e8216558d2afa034516018346060183472601834436012205558dc207e204c58f5d8d83465601834746018344660103447601a206dd8ec2046204458cc18e8216558d2af603459600834686008347a6008344b6002205558dc207e204c58f5d8d8346d6008347c6008344e6000344f600a206dd8ec2046204458cc18e8216558d2af2034516008346060083472600834436002205558dc207e204c58f5d8d83465600834746008344660003467600a206dd8ec2046206458e558e0216518d2aee01551306710b9306711315c18347060083c40600fd167d160505e38897fe33b59700aa9363f597005a863a8b11a03a8613956800629583469501034785018347a5018344b501a206d98ec207e204c58fdd8e0347d5018347c5018344e5010344f50122075d8fc2046204458c418f0217d98e36f983461501034705018347250183443501a206d98ec207e204c58fdd8e0347550183474501834465010344750122075d8fc2046204458c418f0217d98e36f583469500034785008347a5008344b500a206d98ec207e2040347d5000344c500c58fd58f2207418f8344e5000344f50093166600e296c2046204458c418f02175d8f3af10347150083470500834425000344350022075d8fc2046204458c418f83475500834445000344650003457500a207c58f42046205418d5d8d0215598d2aed03c5960103c7860183c7a60183c4b6012205598dc207e204c58f5d8d03c7d60183c7c60183c4e60103c4f60122075d8fc2046204458c418f0217598d2afa03c5160103c7060183c7260183c436012205598dc207e204c58f5d8d03c7560183c7460183c4660103c4760122075d8fc2046204458c418f0217598d2af603c5960003c7860083c7a60083c4b6002205598dc207e204c58f5d8d03c7d60083c7c60083c4e60003c4f60022075d8fc2046204458c418f0217598d2af203c5160003c7060083c7260083c436002205598dc207e204c58f5d8d03c7560083c7460083c4660083c6760022075d8fc204e206c58ed98e8216558d2aee01559306710b130771130dc183c70600834407007d17fd160505e38897fe63e39700b28833b59700aa93468613156600629583469501034785018347a5018344b501a206d98ec207e204c58fdd8e0347d5018347c5018344e5010344f50122075d8fc2046204458c418f0217d98e36f983461501034705018347250183443501a206d98ec207e204c58fdd8e0347550183474501834465010344750122075d8fc2046204458c418f0217d98e36f583469500034785008347a5008344b500a206d98ec207e2040347d5000344c500c58fd58f2207418f8344e5000344f50093166b00e296c2046204458c418f02175d8f3af10347150083470500834425000344350022075d8fc2046204458c418f83475500834445000344650003457500a207c58f42046205418d5d8d0215598d2aed03c5960103c7860183c7a60183c4b6012205598dc207e204c58f5d8d03c7d60183c7c60183c4e60103c4f60122075d8fc2046204458c418f0217598d2afa03c5160103c7060183c7260183c436012205598dc207e204c58f5d8d03c7560183c7460183c4660103c4760122075d8fc2046204458c418f0217598d2af603c5960003c7860083c7a60083c4b6002205598dc207e204c58f5d8d03c7d60083c7c60083c4e60003c4f60022075d8fc2046204458c418f0217598d2af203c5160003c7060083c7260083c436002205598dc207e204c58f5d8d03c7560083c7460083c4660083c6760022075d8fc204e206c58ed98e8216558d2aee01559306710b130771130dc183c70600834407007d17fd160505e38897fe63f797002d4563f4a356850311a0328b13b513003375a8006319055a13146b00638f095ae3765b63b3048c0003c5990183c5890103c6a90183c6b90122054d8d4206e206558e518d83c5d90103c6c90183c6e90103c7f901a205d18dc2066207d98ed58d82154d8d2af903c5190183c5090103c6290183c6390122054d8d4206e206558e518d83c5590103c6490183c6690103c77901a205d18dc2066207d98ed58d82154d8d2af503c5990083c5890003c6a90083c6b90022054d8d4206e206558e518d83c5d90003c6c90083c6e90003c7f900a205d18dc2066207d98ed58d82154d8d2af103c5190083c5090003c6290083c6390022054d8d4206e206558e518d83c5590003c6490083c6690003c77900a205d18dc2066207d98ed58d82154d8d2aed03c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8d2afa03c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8d2af603c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8d2af203c5140083c5040003c6240083c6340022054d8d4206e206558e518d83c5540003c6440083c6640003c77400a205d18dc2066207d98ed58d82154d8d2aee01559305710b1306711301cd83c60500034706007d16fd150505e388e6fe63e5e63a4e89280a13060004e28597800000e780e055130600046285a68597900000e780c0992c0a13060004268597800000e780e05393090c04280913060004e28597800000e780a0520144568b1305fbff6370a414130871139308711b93156400ce954a76aa760a77ea6732fb36f73af33eef03c6950183c6850103c7a50183c7b5012206558e4207e2075d8f598e83c6d50103c7c50183c7e50183c4f501a206d98ec207e204c58fdd8e8216558e32fa03c6150183c6050103c7250183c735012206558e4207e2075d8f598e83c6550103c7450183c7650183c47501a206d98ec207e204c58fdd8e8216558e32f603c6950083c6850003c7a50083c7b5002206558e4207e2075d8f598e83c6d50003c7c50083c7e50083c4f500a206d98ec207e204c58fdd8e8216558e32f203c6150083c6050003c7250083c735002206558e4207e2075d8f598e83c6550003c7450083c7650083c57500a206d98ec207e205dd8dd58d8215d18d2eee81554686c28681cd0347060083c70600fd167d168505e308f7fe6366f7000504e319a4ec2a84637aa4162a8b93146500e2944a75aa750a76ea662afb2ef732f336ef03c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8d2afa03c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8d2af603c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8d2af203c5140083c5040003c6240083c6340022054d8d4206e20683c55400558e498e03c54400a20583c6640003c77400c98d1305fbffc2066207d98ed58d8215d18d2eee81551306711b9306711381cd0347060083c70600fd167d168505e308f7fee365f7ec131a64004e9a280a13060004d28597800000e7802029130600045285a68597800000e780006d2c0a13060004268597800000e78020270504a9b3930414002c0913060004628597800000e780a025e3eb9a10b38a9a409a04269cca8963e47a016fe06f866fe0af80014593d81a0013966a00b304cc00e286130700fcb6873386e4000304060083850700238087002300b6000507850765f70505938404fc93860604e31b15fd134bfbff569b054585b46285d68597200000e78080c40148fd3c6fe0cf816285d68597200000e78040d8e30305a46fd0fffa627c427a11a0568a13097113130d710be3784b076294280a13060004e28597800000e780a01a130600046285a28597800000e780805e2c0a13060004228597800000e780a018930b0c04930afaffa80813060004e28597800000e78020170144131564005e9583459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18d2ef983451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2ef583459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2ef183451500034605008346250003473500a205d18dc2066207d98ed58d034655008346450003476500034575002206558e42076205598d518d02154d8d2aed4675a6750676e6662afa2ef632f236ee01559305710b1306711305c183c60500034706007d16fd150505e388e6fe63f6e6000504e31754ed5684d685ae84637bb41213956400629583459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18d2ef983451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2ef583459500034685008346a5000347b500a205d18dc20662070346d500d98ecd8e8345c50022060347e5008347f5004d8e9385f4ff4207e2075d8f598e0216558e32f1034615008346050003472500834735002206558e4207e2075d8f598e83465500034745008347650003457500a206d98ec20762055d8d558d0215518d2aed46752676867666672afa32f636f23aee01556a86ca86e30105ee0347060083c70600fd167d160505e307f7fee376f7ec63ef845a62fc4ef066e852f863e79a5a814a8149014b814d26e43385844022f493156400de951a05338ca50093030008130300082eecae8b130871079302101033057c41135e650063775e0233b56d01b3b55901c98d3305b040137505f872952a8663e46d011e862a83b28389e513531500b303654063856d01639e5929a1aa630503148145130b81095e859308711b03469501834685010347a5018347b5012206558e4207e2075d8f598e8346d5010347c5018347e5010344f501a206d98ec2076204c18fdd8e8216558e32fb034615018346050103472501834735012206558e4207e2075d8f598e83465501034745018347650103447501a206d98ec2076204c18fdd8e8216558e32f703469500834685000347a5008347b5002206558e4207e2075d8f598e8346d5000347c5008347e5000344f500a206d98ec2076204c18fdd8e8216558e32f3034615008346050003472500834735002206558e4207e20783465500034445005d8f598ea206c18e03476500834775002300bb0085054207e2075d8fd98e8216558e32ef0156c686428715c283c7060003440700b3b48700a18f3334f000b3079040c18f7d17fd160506e5d311a0814713b6f7ff329b13050504e39665ec19a0130b8109930d810963925915638c03120145930a8111e2859308711b2380aa00050503c695fd83c685fd03c7a5fd83c7b5fd2206558e4207e2075d8f598e83c6d5fd03c7c5fd83c7e5fd83c4f5fda206d98ec207e204c58fdd8e8216558e32fb03c615fd83c605fd03c725fd83c735fd2206558e4207e2075d8f598e83c655fd03c745fd83c765fd83c475fda206d98ec207e204c58fdd8e8216558e32f703c695fc83c685fc03c7a5fc83c7b5fc2206558e4207e2075d8f598e83c6d5fc03c7c5fc83c7e5fc83c4f5fca206d98ec207e204c58fdd8e8216558e32f303c615fc83c605fc03c725fc83c735fc2206558e4207e2075d8f598e83c645fc03c755fc83c765fc83c475fc938505fc2207d98ec207e204c58fdd8e8216558e32ef0156c686428701ce83c70600034407007d17fd160506e38887fe33b68700b29ae31f75ec19a0930a8111930981113309bb4133853a416363a9002a896309090cf2e09ee49ae803c50d001a05b385ab00280b1306000497800000e78080bb03ca090003c50d00934cfaff93956c00e2951a05de845e951306000497800000e78040b905456315a900ce8b6e8d99a87d1903c51d00138d1d001a053384a4001345faff136505f01a05629513060004a28597800000e780e0b503ca1900938b1900934cfaff93956c00e29513060004228597800000e780e0b37d19ea8dde89e31909fa13956c0062952c0b1306000497800000e78000b2930d1d0093891b001308710793021010a68b4663a663066e33c56d013335a0007d15337565001a05aa9b33c559013335a000b30570407d156d8d1a052a9ce3725ec263f86d0562840345fbff1309fbff1a05b384ab00130404fc280b13060004a68597800000e78060ab130600042685a28597800000e78040ef2c0b13060004228597800000e78060a94a8be3ee2dfb91a85e8463f8590503c5faff1389faff1345f5ff1a05b304ac00280b13060004a28597800000e78060a6130600042285a68597800000e78040ea2c0b13060004268597800000e78060a413040404ca8ae3ec29fb62653305a4401981a27aaa9aac08130600046274228597800000e780e0a1c27463f99a0c139c6a00229c280a13060004a28597800000e78020a0130600042285e28597800000e78000e42c0a13060004628597800000e780209e33845441568963e38a0022897d1493090c04d54bc26c930d711363fe8a006275d6850276e68697d0ffffe780a07462f0a28a4e8c11a84e85a2856286e68697d0ffffe7802073627c2275a2653335b50013451500aae813d534003335a900134d150056f862fc827963e47a016fd02ff96fd08ff36285d68597100000e780609d6fd0cff35a85d68597a0ffffe780807900005a85d285cdbf5685a685f5b72685ddb72285ddbf5d7186e4a2e026fc8505a5c12a8408659314150063e39500ae84914563e3950091449795000083b5e5fbb3b5b400930640063386d402860509c918603305d5023af0894636f42af811a002f42800141097b0ffffe78020a1a265426581cdfd55fe158505630ab50009ed9760ffffe780a09f000008e004e4a6600664e274616182809760ffffe780809d0000130101dc233c1122233881222334912223302123233c312123384121368483c60600ba84b2892e8a2a89e5ce83c5040085e1138514009705ffff938505dd1306000297800000e780e0c80125630905140a8597200000e78060ad0545230ca1100a852c0a05469760ffffe780801d230c41110a852c0a05469760ffffe780601c0a8513060002ce859760ffffe780601b280aa28597000000e78080130a852c0a130600029760ffffe780a019280aa68597000000e780c0110a852c0a130600029760ffffe780e017280a8a851306800f97700000e780807d1304190002ea02e602e282fd280aac199780ffffe78000d2ac1913060002228597700000e780007b230009008330812303340123833481220339012283398121033a0121130101248280130514009705ffff938505ce1306000297800000e780e0b983c5040001253366b50029e6138514009705ffff9385c5cb1306000297800000e780a0b701250de9130610024a8581458330812303340123833481220339012283398121033a0121130101241773000067004365e31105ea05474a85d2854e86a68631a04a85d2854e86a28601478330812303340123833481220339012283398121033a012113010124170300006700e30f130101dc233c1122233881222334912223302123233c3121ae8483c505002a89d5c51384240093892402280097200000e780009309452300a11228000c1205469760ffffe7802003280013060002a2859760ffffe7802002280013060002ce859760ffffe7802001038514002300a11228000c1205469760ffffe780c0ff08122c001306800f97700000e780606502ee02ea02e602e208120c029780ffffe78020ba0c02130600024a8597700000e7802063833081230334012383348122033901228339812113010124828093851400130600024a85833081230334012383348122033901228339812113010124177300006700e35e130101da233c1124233881242334912423302125233c312323384123b68483c606002e892a84638a061403c5b40383c5a40303c6c40383c6d40322054d8d4206e206558e518d83c5f40303c6e40383c6040483c71404a205d18dc206e207dd8ed58d82154d8daaea03c5340383c5240303c6440383c6540322054d8d4206e206558e518d83c5740303c6640383c6840383c79403a205d18dc206e207dd8ed58d82154d8daae603c5b40283c5a40203c6c40283c6d40222054d8d4206e206558e518d83c5f40203c6e40283c6040383c71403a205d18dc206e207dd8ed58d82154d8daae203c5340283c5240203c6440283c6540222054d8d4206e20683c57402558e518d03c66402a20583c6840283c794024d8e93852400c206e207dd8e558e0216518d2afe05c3131589036d91301a329503060500937679000547b316d700558e2300c500130524001306000297700000e7808049130524022c1a1306000297700000e7806048038514000525a300a40005452300a4007da8b289850402ec02e802e402e005c3131589036d918a852e95830505001376790085463396c600d18d2300b500130a2400081097100000e780a06b230c211308102c1a054605499760ffffe780c0db081013060002ce859760ffffe780c0da081013060002a6859760ffffe780c0d9281a0c101306800f97700000e780603f02fa02f602f202ee281a2c0a9780ffffe78020942c0a13060002528597700000e780203d130524028a851306000297700000e780003ca3002401230024018330812503340125833481240339012483398123033a0123130101268280157186eda2e9a6e5cae14efd52f956f55af15eed62e966e5328a7d16637ab63c2e89637aba3aaa89930a7102130b7108930b7108130c71065284050a93146400ce9403c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8d2ae103c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8daafc03c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8daaf803c5140083c5040003c6240083c6340022054d8d4206e206558e518d83c5540003c6440083c6640003c77400a205d18dc2066207d98ed58d82154d8daaf403c594fd83c584fd03c6a4fd83c6b4fd22054d8d4206e206558e518d83c5d4fd03c6c4fd83c6e4fd03c7f4fda205d18dc2066207d98ed58d82154d8d2af003c514fd83c504fd03c624fd83c634fd22054d8d4206e206558e518d83c554fd03c644fd83c664fd03c774fda205d18dc2066207d98ed58d82154d8d2aec03c594fc83c584fc03c6a4fc83c6b4fc22054d8d4206e206558e518d83c5d4fc03c6c4fc83c6e4fc03c7f4fca205d18dc2066207d98ed58d82154d8d2ae803c514fc83c504fc03c624fc83c634fc22054d8d4206e20683c554fc558e518d03c644fca20583c664fc03c774fcd18d938c04fcc2066207d98ed58d82154d8d2ae40155da855686630b051883c60500034706007d16fd150505e387e6fe63f0e618280013060004a68597700000e7804013130600042685e68597700000e78040127d14630504147d1493146400ce940275e2654266a266aaf0aeecb2e8b6e403c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8d2ae103c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8daafc03c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8daaf803c5140083c5040003c6240083c6340022054d8d4206e206558e518d83c5540003c6440083c6640003c77400a205d18dc2066207d98ed58d82154d8daaf40155e2855e8605c983c60500034706007d16fd150505e388e6fe63fee600130600046685a68597700000e78000fea68ce31004ecce8c2c0013060004668597700000e78080fce3132ac7ee604e64ae640e69ea794a7aaa7a0a7bea6b4a6caa6c2d61828017f5feff1305e5569305e0029790ffffe78060540000317106fd22f926f54af14eed52e956e55ae1defce2f8e6f4eaf02e89aa8993da1500130bf103930bf101130cf103930cf101fd1a13961a00130816006377284956850906637f262193166800ce9603c7960183c7860183c4a60103c4b60122075d8fc2046204458c418f83c7d60183c4c60103c4e60183c5f601a207c58f4204e205c18ddd8d8215d98d2eec83c5160103c7060183c7260183c43601a205d98dc207e204c58fdd8d03c7560183c7460183c4660103c4760122075d8fc2046204458c418f0217d98d2ee883c5960003c7860083c7a60083c4b600a205d98dc207e20403c7d60003c4c600c58fdd8d2207418f83c7e60083c4f6001a064e96c207e204c58f5d8f0217d98d2ee483c5160003c7060083c7260083c43600a205d98dc207e204c58fdd8d03c7560083c7460083c4660083c6760022075d8fc204e206c58ed98e8216d58d2ee083459601834686010347a6018347b601a205d58d4207e2075d8fd98d8346d6010347c6018347e6018344f601a206d98ec207e204c58fdd8e8216d58d2efc83451601834606010347260183473601a205d58d4207e2075d8fd98d83465601034746018347660183447601a206d98ec207e204c58fdd8e8216d58d2ef883459600834686000347a6008347b600a205d58d4207e2075d8fd98d8346d6000347c6008347e6008344f600a206d98ec207e204c58fdd8e8216d58d2ef483451600834606000347260083473600a205d58d4207e2075d8fd98d83465600034746008347660003467600a206d98ec20762065d8e558e0216d18d2ef00156de865a8719ce83c70600834407007d17fd160506e38897fe33ba970021a0428a19a0014a429a6379257763742a771a053384a90093146a00ce9403459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8d2aec0345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8d2ae803459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8d2ae40345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8d2ae003c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8d2afc03c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8d2af803c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8d2af403c5140083c5040003c6240083c6340022054d8d4206e206558e518d83c5540003c6440083c6640003c77400a205d18dc2066207d98ed58d82154d8d2af00155e685628639c983c60500034706007d16fd150505e388e6fe63f1e604081013060004a28597700000e78080af130600042285a68597700000e78060f30c1013060004268597700000e78080ad13161a00130816005285e36e28b7e3940ab6130bf103930bf101130cf103930cf101094dca8afd1a63fb2a4f13946a004e94081013060004ce8597700000e78060a9130600044e85a28597700000e78040ed0c1013060004228597700000e78060a763ebaa490146014505480906637f562193166800ce9603c7960183c7860183c4a60103c4b60122075d8fc2046204458c418f83c7d60183c4c60103c4e60183c5f601a207c58f4204e205c18ddd8d8215d98d2eec83c5160103c7060183c7260183c43601a205d98dc207e204c58fdd8d03c7560183c7460183c4660103c4760122075d8fc2046204458c418f0217d98d2ee883c5960003c7860083c7a60083c4b600a205d98dc207e20403c7d60003c4c600c58fdd8d2207418f83c7e60083c4f6001a064e96c207e204c58f5d8f0217d98d2ee483c5160003c7060083c7260083c43600a205d98dc207e204c58fdd8d03c7560083c7460083c4660083c6760022075d8fc204e206c58ed98e8216d58d2ee083459601834686010347a6018347b601a205d58d4207e2075d8fd98d8346d6010347c6018347e6018344f601a206d98ec207e204c58fdd8e8216d58d2efc83451601834606010347260183473601a205d58d4207e2075d8fd98d83465601034746018347660183447601a206d98ec207e204c58fdd8e8216d58d2ef883459600834686000347a6008347b600a205d58d4207e2075d8fd98d8346d6000347c6008347e6008344f600a206d98ec207e204c58fdd8e8216d58d2ef483451600834606000347260083473600a205d58d4207e2075d8fd98d83465600034746008347660003467600a206d98ec20762065d8e558e0216d18d2ef00156de865a8719ce83c70600834407007d17fd160506e38897fe33ba970021a0428a19a0014a429a63715529637e5a271a053384a90093146a00ce9403459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8d2aec0345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8d2ae803459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8d2ae40345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8d2ae003c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8d2afc03c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8d2af803c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8d2af403c5140083c5040003c6240083c6340022054d8d4206e206558e518d83c5540003c6440083c6640003c77400a205d18dc2066207d98ed58d82154d8d2af00155e6856286e30405b883c60500034706007d16fd150505e387e6fee3f9e6b6081013060004a28597600000e7800061130600042285a68597700000e780e0a40c1013060004268597600000e780005f13161a00130816005285e36d58b705beea704a74aa740a79ea694a6aaa6a0a6be67b467ca67c067d296182805285d68529a0528511a05685ca859790ffffe780403f0000757106e522e1a6fccaf8cef4d2f0d6ecdae8dee4ae89fd1513d61500d18d13d62500d18d13d64500d18d13d68500d18d13d60501d18d13d60502d18d93c5f5ff17860000033686c19786000083b686c113d71500798e918d33f6d5008981f58db29517860000033666c09786000083b666c013d74500ba95f18db385d502e1917d56b35ab600850a638a0a0a2a8913d519007999fd1a130bf5ff13d529001e054a95130405fc8d44ce8b63723b091395db0033457501935575002d8d93151501b3cba50033f55b01b3353501fd15b3f535010d8d637e35051a05330aa900280013060004a28597600000e780e04b130600042285d28597700000e780c08f2c0013060004528597600000e780e049050bfd1413040404d1f8aa600a64e6744679a679067ae66a466ba66b496182805a85ce859790ffffe780802b000017f5feff130545a1f1459790ffffe780e0a00000557186e5a2e126fd4af94ef552f156ed5ae95ee562e1e6fceaf8eef42e8c2a89014b930b7104930c710213bd2503954d854463f384238545139564004a9503469501834685010347a5018347b5012206558e4207e2075d8f598e8346d5010347c5018347e5010344f501a206d98ec2076204c18fdd8e8216558e32f0034615018346050103472501834735012206558e4207e2075d8f598e83465501034745018347650103447501a206d98ec2076204c18fdd8e8216558e32ec03469500834685000347a5008347b5002206558e4207e2075d8f598e8346d5000347c5008347e5000344f500a206d98ec2076204c18fdd8e8216558e32e8034615008346050003472500834735002206558e4207e2075d8f598e83465500034745008347650003447500a206d98ec2076204c18fdd8e8216558e32e4034695fd834685fd0347a5fd8347b5fd2206558e4207e2075d8f598e8346d5fd0347c5fd8347e5fd0344f5fda206d98ec2076204c18fdd8e8216558eb2e0034615fd834605fd034725fd834735fd2206558e4207e2075d8f598e834655fd034745fd834765fd034475fda206d98ec2076204c18fdd8e8216558e32fc034695fc834685fc0347a5fc8347b5fc2206558e4207e2075d8f598e8346d5fc0347c5fc8347e5fc0344f5fca206d98ec2076204c18fdd8e8216558e32f8034615fc834605fc034725fc834735fc2206558e4207e2075d8f598e834655fc034745fc834765fc034575fca206d98ec20762055d8d558d0215518d2af401556686de8601cd0347060083c70600fd167d160505e308f7fe6369f7008504b3b58401e39384df51a0814533c58401133515003366ad003dea9389f4ff63f789098589d1c5139a69004a9a939a6400ca9a281013060004d28597600000e780c01c130600045285d68597600000e780c01b2c1013060004568597600000e780c01a0545637f95004a85a6854e8697f0ffffe78060e04a85a68597000000e7804004050be310bbd7014511a00545ae600e64ea744a79aa790a7aea6a4a6baa6b0a6ce67c467da67d696182804e8511a02685e2859790ffffe78080f90000317106fd22f926f54af14eed52e956e55ae12e89aa840345950583c5840503c6a40583c6b40522054d8d4206e206558e518d83c5d40503c6c40583c6e40503c7f405a205d18dc2066207d98ed58d82154d8daafc03c5140583c5040503c6240583c6340522054d8d4206e206558e518d83c5540503c6440583c6640503c77405a205d18dc2066207d98ed58d82154d8daaf803c5940483c5840403c6a40483c6b40422054d8d4206e206558e518d83c5d40403c6c40483c6e40403c7f404a205d18dc2066207d98ed58d82154d8daaf403c5140483c5040403c6240483c6340422054d8d4206e206558e518d83c5540403c6440483c6640403c77404a205d18dc2066207d98ed58d82154d8daaf003c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8d2aec03c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8d2ae803c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8d2ae403c5140083c5040003c6240083c6340022054d8d4206e20683c55400558e518d03c64400a20583c6640003c77400d18d93890404c2066207d98ed58d82154d8d2ae01305f10181551306f1076380051a83460600034705007d157d168505e387e6fe63f5e6180a8513060004a68597600000e78020f1130600042685ce8597600000e78020f00d45636aa914130af107894a130bf10513946a00269403459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8daaec0345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8daae803459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8daae40345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8daae06265c26522668266aafcaef8b2f4b6f00155da8552860dc983c60500034706007d16fd150505e388e6fe63ffe600850a130504fc13060004a28597600000e78020dba289e39f2aeb8a85130600044e8597600000e780c0d9ea704a74aa740a79ea694a6aaa6a0a6b29618280257106ef22eb26e74ae32a8484004800130901031306c002814597600000e78080c9130680132685814597600000e78080c817e5feff9305350441464a8597600000e78020d4370501011b0505022ac082fe8a8522859740ffffe780a056fa605a64ba641a691d6182805d7186e4a2e026fc8505a5c12a8408659314150063e39500ae84914563e3950091449775000083b5853cb3b5b400930600053386d4028e0509c918603305d5023af0a14636f42af811a002f4280014109790ffffe78040dfa265426581cdfd55fe158505630ab50009ed9740ffffe780c0dd000008e004e4a6600664e274616182809740ffffe780a0db00005d7186e4a2e026fc4af8ae84806590612a892800a2859780ffffe780808a0345810001c9426505c59780ffffe780e0b0000005040dc49305910080e4130519001306000297600000e78060c405452300a900a6600664e27442796161828017e5feff1305851df1459780ffffe780201d0000130101d0233c112e2338812e2334912e2330212f233c312d2338412d930700026317f628ba89368a2a8903c5950103c6850183c6a50103c7b5012205518dc2066207d98e558d03c6d50183c6c50103c7e50183c7f5012206558e4207e2075d8f598e0216518d2aec03c5150103c6050183c6250103c735012205518dc2066207d98e558d03c6550183c6450103c7650183c775012206558e4207e2075d8f598e0216518d2ae803c5950003c6850083c6a50003c7b5002205518dc2066207d98e558d03c6d50083c6c50003c7e50083c7f5002206558e4207e2075d8f598e0216518d2ae403c5150003c6050083c6250003c735002205518dc2066207d98e558d03c6550083c6450003c7650083c575002206558e4207e205d98dd18d82154d8d2ae0880a9770ffffe7802041a8088a859770ffffe780e02d766511c556659740ffffe78080be267586756666aae4aee032fc0305711883056118b674034651182303a102a20503452118d18d2312b10283451118220503463118830641184d8d56744206e206558e518d2ad0a808d2854e869770ffffe780c02c11c426859740ffffe78080b86275e6650666aaea26658676b2ee2676aaf2aef6b6fab2fe09452300a118130511180c101d4697600000e780c0a408108c0a9770ffffe780803d880a97000000e780c00e82e882e482e002fc000bc80a04031306c002814597600000e780c094130680132285814597600000e780c09317e5feff930575cf4146268597600000e780609f370501011b0505022328a1142334012ca8088c0a9740ffffe780a02102744276a808a2859740ffffe7800036880aac081306800f97600000e780a09b880a2c189760ffffe780e0f02c18130600024a8597600000e780e099227511c522859740ffffe780e0a98330812f0334012f8334812e0339012e8339812d033a012d13010130828017e5feff130545f697e5feff9386e5fc9305b002900a9780ffffe780400b0000411106e422e02a84086511c508609740ffffe780a0a4087009c9086ca260026441011743ffff670063a3a260026441018280697106f622f226ee4aea4ee652e2d6fddaf9def5e2f1e6ed2e8a2a89014481490d45aae082e49304110501163335c00093b51500b36ab500130b1108894b7d5c88088c009790ffffe7800054034501056309751f6301051003c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8d2ae903c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8d2ae503c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8d2ae103c5140083c5040003c6240083c6340022054d8d4206e206558e518d83c5540003c6440083c6640003c77400a205d18dc2066207d98ed58d82154d8daafc63890a00dda002e902e502e182fc639e0a0ca81813060002d28597600000e78060bd012579e1639a091628110d46a2859770ffffe780804c2a7559c96a75ca752a76aae9aee5b2e1a8188c019790ffffe78000250305eb008305db000346cb00e6792303a10aa205d18d2312b10a03459b0083458b000346ab008306bb0022054d8d4206e206558e518d2ad103451b0083450b0003462b0083463b0022054d8d4206e20683455b00558e518d03464b00a20583466b0003477b00d18d834c0108c2066207d98ed58d82154d8d2aed11a081496a658a550316410a8306610a2af82edc231ec102230fd102630e8409050401b5638609060305e1038315c1036256c2762307a1022316b10232d436f0130511010c103d4697500000e780206b4ee423089101a8182c0005469790ffffe78060d9667535c92a658a656676aaf0aeecb2e888089790ffffe78060f42334a9004e859790ffffe78040a7014531a01305a005a300a90005452300a900b2701274f2645269b269126aee7a4e7bae7b0e7cee6c5561828017e5feff1305e5bef1459780ffffe78080be000017e5feff1305a5f19305b002edb717e5feff1305a5c197d5feff938645489305b00290089780ffffe780a0d60000497186f6a2f2a6eecaeacee6d2e256fe5afa5ef662f266ee6aea6ee62e842ae0814a014d0149014b0945aaf882fc93041108bd497d5a2ee408018c1897000000e780a09303450108630b052803c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8daae103c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8d2afd03c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8d2af903c5140083c5040003c6240083c6340022054d8d4206e206558e518d83c5540003c6440083c6640003c77400a205d18dc2066207d98ed58d82154d8d2af5281113060002a28597600000e780c08d01256310051888190946d6859770ffffe780001dce7b638a0b1e126c6e7563fc8915aae8eaec414581459780ffffe78080672a842e8b4146de8597500000e780204783458400834994000349a400834db4000346c400034dd4008347e400034af400834c04000347140083432400834634000348440003435400834864008342740063050b04228542f0468416fc6aec1a8d4ae81e896ef4b68dcee0ba89b2e452f83e8a2e8b9730ffffe7804051da85d287427a26664e878669ee86a27dca8342696a83626de272a28802786665631e0514a20933e5b9004209e20db3e52d014d8d220db365cd0013960701620a3366ca00d18d8215b3eda50013158700336595019395030113968601d18d4d8d93158300b3e505011396080193968201558ed18d8215b3eca50013040cff93890b01228581459780ffffe780e0562a8c2e8bce85228697500000e7808036e2f9dafd22e2a8098c199790ffffe780a0e28c1188618c65014b6e6daaf0aef405492264bd497d5a466511c55e859730ffffe7800044638a4a07850ab1bb3365690119cd630d0d0226758675026608f20cee233096012334b6012338a6013da01305500382652380a50023b80500630f0d006a859780ffffe780a06e01a81305200382652380a50023b80500b6701674f6645669b669166af27a527bb27b127cf26c526db26d7561828017e5feff13052586f1459780ffffe780c085000017e5feff1305c58997e5feff9386658c9305b002b0099780ffffe780c09e000017e5feff130595b993059002e9b7097186fea2faa6f6caf2ceeed2ead6e6dae25efe62fa66f66af26eeeb289ae842ae4014b014d0149814b32e102e5130411093d4afd5a32ec2ee808090c0197f0ffffe780c05a03450109630c052803459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8daae90345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8daae503459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8daae10345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8d2afd281913060002a68597500000e780e0540125631105180802da854e869770ffffe78020e4126c630b0c1ed26c3265637d9a15aaf0eaf4414581459780ffffe780a02eaa84ae8b4146e28597500000e780400e83c5840003ca940003c9a40083c9b40003c6c40083cdd40083c7e40083caf40003cd040003c7140083c3240083c6340003c8440003c3540083c8640083c2740063850b042685c28bc684d6e016f86ef49a8d4af01e89b6e4d2e83a8ab2ec4efcbe89ae8a9730ffffe7806018d685ce87e27966665287466aa666ca8302796e83a27dc272866aa6885e882675631f0514220a3365ba004209e209b3e529014d8da20db3e5cd0013960701e20a33e6ca00d18d82154d8daaf4131587003365a5019395030113968601d18d4d8d93158300b3e505011396080193968201558ed18d8215b3eda50093840cff130a0c01268581459780ffffe780001eaa8cae8bd285268697500000e780a0fd66e25ee626eaa8110c029790ffffe780c0a98c1988618c65814b2e7daaf8aefc0549e269c2643d4afd5a067511c562859730ffffe780000b630a5b07050ba9bb3365790119cd630d0d026675c675226608f20cee2330b601267508e62338a6013da013055003a2652380a50023b80500630f0d006a859780ffffe780a03501a813052003a2652380a50023b80500f6705674b6741679f669566ab66a166bf27b527cb27c127df26d1961828017d5feff1305254df1459770ffffe780c04c000017d5feff1305c55097d5feff938665539305b002b0119770ffffe780c065000017e5feff130525839305c002e9b7097186fea2faa6f6caf2ceeed2ead6e6dae25efe62fa66f66af26eeeae892ae4014b814a214a52e802ec02f005452af402f8130d9103930d110b0944fd5428182c109790ffffe780e0b0034581036309853475cd03459d0183458d010346ad018346bd0122054d8d4206e206558e518d8345dd010346cd018346ed010347fd01a205d18dc2066207d98ed58d82154d8daae503451d0183450d0103462d0183463d0122054d8d4206e206558e518d83455d0103464d0183466d0103477d01a205d18dc2066207d98ed58d82154d8daae103459d0083458d000346ad008346bd0022054d8d4206e206558e518d8345dd000346cd008346ed000347fd00a205d18dc2066207d98ed58d82154d8d2afd03451d0083450d0003462d0083463d0022054d8d4206e206558e518d83455d0003464d0083466d0003477d00a205d18dc2066207d98ed58d82154d8d2af929a082e582e102fd02f9081913060002ce8597500000e780e01a01256318052208190546da859770ffffe780609a0345010b6311052603c59d0183c58d0103c6ad0183c6bd0122054d8d4206e206558e518d83c5dd0103c6cd0183c6ed0103c7fd01a205d18dc2066207d98ed58d82154d8daafc03c51d0183c50d0103c62d0183c63d0122054d8d4206e206558e518d83c55d0103c64d0183c66d0103c77d01a205d18dc2066207d98ed58d82154d8daaf803c59d0083c58d0003c6ad0083c6bd0022054d8d4206e206558e518d83c5dd0003c6cd0083c6ed0003c7fd00a205d18dc2066207d98ed58d82154d8daaf403c51d0083c50d0003c62d0083c63d0022054d8d4206e206558e518d83c55d0003c64d0083c66d0003c77d00a205d18dc2066207d98ed58d82154d8daaf008190546da859770ffffe7804099ca7b63870b168e653d456378b51a6a79138405ff138c0b01228581459780ffffe78060e3aa84ae8ce285228697500000e78000c326f966fda2e108010c199780ffffe780206f28090c019730ffffe780c01008020c010d469780ffffe780c02f1265630305125265b2651266aae12efd32f908020c199780ffffe780e0595265d145631cb510126451468809a28597500000e780e0bc3265fd5411c522859730ffffe780c0cc0675a67546762af92efdb2e16675aa750a76ea666267aae5a8110ce910e514e1639aea000808d68597f0ffffe78080e7827a426a0944130500053385aa0252950c191306000597500000e78000b70a65850a56f09780ffffe78000f6630709005e859730ffffe78020c6630a9b02050b45b10275e2654266a26688ea8ce690e2f6705674b6741679f669566ab66a166bf27b527cb27c127df26d1961828017d5feff1305450cf1459770ffffe780e00b000017d5feff1305e50f97d5feff938685129305b002901089a017d5feff1305650e97d5feff938605119305b00210022da017d5feff1305e50c97d5feff9386859309a817d5feff1305c50b97d5feff938665129305b00210199770ffffe780c020000041459780ffffe780608e0000757106e522e1a6fccaf8cef4d2f02a89814432e402e81304910181153335b00093351900b369b500094a28082c009780ffffe780406d0345810165d9630c451303459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8daaec0345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8daae803459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8daae40345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8daae0e39909ee880013060002ca8597500000e780a0d70125e31e05ec93f4f40f850413f5f40fe30795ec17d5feff130525eef1459770ffffe780c0ed00002685aa600a64e6744679a679067a49618280517186f5a2f1a6edcae9cee5d2e156fd5af95ef562f166ed6ae96ee5b2892e8a2ae0014b814a32ec02f013049102894d7d5928102c089780ffffe7806054034581026300b51b75cd03459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8daaf40345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8daaf003459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8daaec0345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8daae829a082f482f082ec82e8880813060002d28597500000e78060be012519c1d684a5a88808da854e869760ffffe780804dc66b63820b0c666d8674268581459780ffffe7808098aa8c2e8cde85268697400000e7802078e6e8e2eca6f088188c089780ffffe7804024ac1888618c65c674aae8aeec63870a0056859780ffffe78040b56665c6652ae82ee463070d005e859730ffffe780e08463052b05050ba68a89bd63890a004265a265026608ea32850ce639a01305b00682652384a5002e8523305501ae700e74ee644e69ae690e6aea7a4a7baa7b0a7cea6c4a6daa6d6d61828017d5feff1305a5c9f1459770ffffe78040c9000017d5feff130545cd97d5feff9386e5cf9305b00290189770ffffe78040e20000357106ed22e926e5aa85a8100d4697000000e780c0d9267461c88304010793051107130511013d4697400000e780206922e423089100a8102c0011469780ffffe78060d726754dcd6675c67526762af82ef432f0a8100c1001469780ffffe78080d526755dc56675c6752676aae4aee032fc88082c1809469780ffffe780a0d3466545c50675e6654666aafcaef8b2f4231201088808ac105001894689449780ffffe78000a70345010541ed6665631b950a8314410826759780ffffe78000a062759780ffffe780609f02759780ffffe780c09e22859780ffffe780209e014501469b95040131a003450107814522050546d18d4d8dea604a64aa640d61828017d5feff130545bb97c5feff9386e54109a817d5feff130525ba97c5feff9386c5409305b00290080da817d5feff1305a5b897c5feff9386453f9305b002b01029a817d5feff130525b797d5feff9386458e9305b002130671089770ffffe78000cc000017d5feff130585a0b9459770ffffe780c0af0000517186f5a2f1a6edcae9cee5d2e156fd5af95ef562f166ed6ae96ee5b2892e8a2ae0014b814a32ec02f013049102894d7d5928102c089780ffffe7808017034581026300b51b75cd03459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8daaf40345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8daaf003459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8daaec0345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8daae829a082f482f082ec82e8880813060002d28597500000e7808081012519c1d684a5a88808da854e869760ffffe780a010c66b638a0b0a666d8674268581459770ffffe780a05baa8c2e8cde85268697400000e780403be6e8e2eca6f088188c089780ffffe78060e7ac1888618c65c674aae8aeec63870a0056859770ffffe78060786665c6652ae82ee463070d005e859720ffffe7800048630d2b03050ba68a89bd63820a064265a265026608ea0ce623305601ae700e74ee644e69ae690e6aea7a4a7baa7b0a7cea6c4a6daa6d6d61828017d5feff1305c58df1459770ffffe780608d000017d5feff1305659197d5feff938605949305b00290189770ffffe78060a6000017d5feff1305a5879305b002e9b7130101ce233c1130233881302334913023302131233c312f2338412f2334512f2330612f233c712d2338812d2334912d2330a12d233cb12b3a8a3684328bae892a891305000285459720ffffe780c03a6306056eaa8413060002814597400000e780401c514585459720ffffe780c0386306056c2a8c5146814597400000e780601a1305000281459770ffffe780c045aa8bae8a13060002d28597400000e780402526859720ffffe78080350345140183450401034624018306340122054d8d4206e206558e518daac803459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8daae40345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8daae0130a0105930c8104514581459770ffffe78020392afeaee282e693041104281a8c0026869770ffffe780401e13042104281aa68522869770ffffe780201d93043104281aa28526869770ffffe780001cc000281aa68522869770ffffe780001b93045104281aa28526869770ffffe780e01913046104281aa68522869770ffffe780c01893047104281aa28526869770ffffe780a017281aa68566869770ffffe780c01613049104281ae68522869770ffffe780a0159304a104281aa28526869770ffffe78080141304b104281aa68522869770ffffe7806013e400281aa28526869770ffffe78060121304d104281aa68522869770ffffe78040119304e104281aa28526869770ffffe78020101304f104281aa68522869770ffffe780000f281aa28552869770ffffe780200e13041105281ad28522869770ffffe780000d93042105281aa28526869770ffffe780e00b13043105281aa68522869770ffffe780c00ad008281aa2859770ffffe780e009f27c966d366a62859720ffffe780c0131304ca02636e4445228581459770ffffe78000212afeaee282e64145a1459720ffffe780e010630705442a8c31452330ac001305c0022334ac00a2c0d000281a8c009770ffffe78040048944130d410462840860aac0281a8c006a869770ffffe780a002fd142104edf462859720ffffe780800c13860b02281ade859770ffffe780a00033864c01281ae6859770ffffe780a0ff727a166d366c63870a005e859720ffffe780400963870d0066859720ffffe78060085a8581459770ffffe78020162a84ae8ace855a8697400000e780c0f5130500026314ab3a03056400230fa112030554008345440022054d8d231ea1120345140083450400034624008306340022054d8d4206e206558e518d232ca1120345840083457400034694008346a40022054d8d4206e206558e518d8345c4000346b4008346d4000347e400a205d18dc2066207d98ed58d8215b3e9a500034504018345f400034614018346240122054d8d4206e206558e518d83454401034634018346540103476401a205d18dc2066207d98ed58d8215b3eba5000345840183457401034694018346a40122054d8d4206e206558e518d8345c4010346b4018346d4010347e401a205d18dc2066207d98e034bf401d58d8215b3e4a50063870a0022859720ffffe780e0f50305e1138315c113032681132303a1042312b104b2c0a303310513d589032307a10413d50903a306a10413d589022306a10413d50902a305a10413d589012305a10413d50901a304a10413d589002304a104a307710513d58b03230ba10413d50b03a30aa10413d58b02230aa10413d50b02a309a10413d58b012309a10413d50b01a308a10413d58b002308a104a30b910413d58403230fa10413d50403a30ea10413d58402230ea10413d50402a30da10413d58401230da10413d50401a30ca104a180230c9104a30f6105281a9750ffffe780806908108c009750ffffe7804056166511c572759720ffffe780e0e64275a27502762aec2ee832e40305f1168305e11656640346d1162303a100a2050345a116d18d2312b1008345911622050346b1168306c1164d8df6644206e206558e518d2ac00810d28562869750ffffe780205591c422859720ffffe780e0e02265827542662afe6265a276b2e24276aae6aeeab6eeb2f205452304a116130591168a851d4697400000e78020cd28002c1a9750ffffe780e065281a97e0ffffe780203702fc02f802f402f0a01a681aa4121306c002814597400000e78020bd130680132285814597400000e78020bc17c5feff9305d5f74146268597400000e780c0c7370501011b050502232ca1122338012a88002c1a9720ffffe780004a226462668800a2859720ffffe780605e281a8c001306800f97400000e78000c4281a0c109740ffffe78040190c10130600024a8597400000e78040c2426511c522859720ffffe78040d263070d0052859720ffffe78060d1833081310334013183348130033901308339812f033a012f833a812e033b012e833b812d033c012d833c812c033d012c833d812b13010132828017c5feff130525a5f1459760ffffe780c01600009720ffffe78080cd000017c5feff1305251a97c5feff9386c51e9305b002301a9760ffffe780202f0000130101dd2334112223308122233c91202e84aa8402f002ec02e802e4281097e0ffffe780a0de22f228100c1221469720ffffe780004f08122c101306800f97400000e780a0b408122c009740ffffe780e0092c0013060002268597400000e780e0b2833081220334012283348121130101238280130101812334117e2330817e233c917c2338217d2334317d2330417d233c517b2338617b2334717b2330817b233c91792338a1792334b179357136ec32e42ee82a842338014623340146a80813068002814597400000e780409f0335014683358146033601472ae12ee5086032e902f10c683336a00014643307c040f98d32f502f92afdb6e1b2e582e9aaedb6f1aef5130da122930ba124854d930a400828119770ffffe780207519e16f2090222a8493040501233c0178233801782334017823300178881697e0ffffe780e0cc88165146a6859720ffffe780603d130501468c161306800f97400000e780e0a213050146930501789740ffffe780e0f7033581798335017903368178833601782ae62ee2b2fdb6f9033b0400033c84002af62ef232ee36ea233c0178233801782334017823300178881697e0ffffe780c0c5233481472330614788169305014641469720ffffe780a035130501468c161306800f97400000e780209b13050146930501789740ffffe78020f0930501781306000213041113228597400000e780c0982308011217c5feff9305e5ed13060002228597400000e780a0d9012521c1327592757266d2664a6a2334a1282330b128233cc1262338d12663080a046a648c1c52859780ffffe780c083ae842dcd41c48e04d29403ba04227d14d5b74a64e30a04386a65b384ad400c0a22859780ffffe780208163000518e38db4378e05a29503b405228504cdb7833981278334012803398128033401279770ffffe780a068233805208545231db52000e12334350104e9233c250123348517233065172ae902ed6f00f0329204d29423b4841723b064176f001032033d812783350128833c81280359aa21833b01272d456379a91293891400139454005294939a44006375391d2300740113d58b03a303a40013d50b032303a40013d58b02a302a40013d50b022302a40013d58b01a301a40013d50b012301a40013d58b00a300a4002304a40113558d03a307a40013550d032307a40013558d02a306a40013550d022306a40013558d01a305a40013550d012305a40013558d00a304a4002308b40013d58503a30ba40013d50503230ba40013d58502a30aa40013d50502230aa40013d58501a309a40013d505012309a40013d58500a308a400230c940113d58c03a30fa40013d50c03230fa40013d58c02a30ea40013d50c02230ea40013d58c01a30da40013d50c01230da40013d58c00a30ca400f5aa2300015a639ab40323308136233401362338b136130501468c161306015a9770ffffe780806d6f20206f854d1545aee463f2a41e1149e5aa8e05a29503b5052299c8b30590400356a5210e06329503350522fd15edf98355a521fd152338a164233c01642330b16613050146930501651306015a9770ffffe78020680335814783350147233ca17803368146833601462338b178033501492334c1782330d1780339014a8355a521833481492a846374b9006f20004e0334052119e06f20204d035985218355a42185042285e375b9fe6f20204c139559005295b304994013965400d6e8ae8aa28597400000e78060af13d58b03a303a40013d50b032303a40013d58b02a302a40013d50b022302a40013d58b01a301a40013d50b012301a40013d58b00a300a4002300740113558d03a307a40013550d032307a40013558d02a306a40013550d022306a40013558d01a305a40013550d012305a40013558d00a304a4002304a40113d58a03a30ba40013d50a03230ba40013d58a02a30aa40013d50a02230aa40013d58a01a309a40013d50a012309a40013d58a00a308a40023085401c66a13d58c03a30fa40013d50c03230fa40013d58c02a30ea40013d50c02230ea40013d58c01a30da40013d50c01230da40013d58c00a30ca400230c940113050a16b305550192094e951396440097400000e780c09e0529d29a23b48a1723b06a17231d2a21130da122930ba124cda76389a400814d19456397a4008144154929a0268919a0e5141949e2e09770ffffe780e02faa8a23380520231d05200355aa219349f9ffaa99239d3a2193155900d29503c6950183c6850103c7a50183c7b5012206558e4207e2075d8f598e83c6d50103c7c50183c7e50103c4f501a206d98ec2076204c18fdd8e8216558e233cc14603c6150183c6050103c7250183c735012206558e4207e2075d8f598e83c6550103c7450183c7650103c47501a206d98ec2076204c18fdd8e8216558e2338c14603c6950083c6850003c7a50083c7b5002206558e4207e2075d8f598e83c6d50003c7c50083c7e50003c4f500a206d98ec2076204c18fdd8e8216558e2334c14603c6150083c6050003c7250083c735002206558e4207e2075d8f598e83c6550003c7450083c7650083c57500a206d98ec207e205dd8dd58d8215d18d2330b146b14563e4b9006f30802dca8613041900018d630435016f30e02c5a8c6689930c0a161395460066950c65aee808612afc93155400d295139659005685368b97300000e780c03f93154400e69513850a161396490097300000e780603e231d6a21033501468335814603360147833681472330a1362334b1362338c136233cd136528663930d0056860357a6219389140013945400329493974400ca8c628b637c370f2300740113d58b03a303a40013d50b032303a40013d58b02a302a40013d50b022302a40013d58b01a301a40013d50b012301a40013d58b00a300a4002304a40113558d03a307a40013550d032307a40013558d02a306a40013550d022306a40013558d01a305a40013550d012305a40013558d00a304a400a6652308b40013d58503a30ba40013d50503230ba40013d58502a30aa40013d50502230aa40013d58501a309a40013d505012309a40013d58500a308a400230c940113d58c03a30fa40013d50c03230fa40013d58c02a30ea40013d50c02230ea40013d58c01a30da40013d50c01230da40013d58c00a30ca40005aa139559003295b30d9740328913965d00a2853a8cbe8497300000e780c06d13d58b03a303a40013d50b032303a40013d58b02a302a40013d50b022302a40013d58b01a301a40013d50b012301a40013d58b00a300a4002300740113558d03a307a40013550d032307a40013558d02a306a40013550d022306a40013558d01a305a40013550d012305a40013558d00a304a4002304a401a66513d58503a30ba40013d50503230ba40013d58502a30aa40013d50502230aa40013d58501a309a40013d505012309a40013d58500a308a4002308b40013d58c03a30fa40013d50c03230fa40013d58c02a30ea40013d50c02230ea40013d58c01a30da40013d50c01230da40013d58c00a30ca400230c940113050916b305950092094e9513964d0097300000e780205da68762874a86c66de27486661b051700b305f60023b4d51623b06517231da62003358137833501370336813683360136233ca1782338b1782334c1782330d178233ca15a2338b15a2334c15a2330d15a03350a216309052c8149d687268c6e8d03598a218335815b0336015b8336815a0337015a233cb1782338c1782334d1782a8a2330e178835ba5212d4563ebab32cee4054b91491545bee0636fa9006309a900014b19456317a9000149954929a0ca8919a0651999499770ffffe78060e8aa8a23380520231d05200355aa2113c4f9ffb30ca400239d9a2193955900d29503c6950183c6850103c7a50183c7b5012206558e4207e2075d8f598e83c6d50103c7c50183c7e50183c4f501a206d98ec207e204c58fdd8e8216558e233cc14603c6150183c6050103c7250183c735012206558e4207e2075d8f598e83c6550103c7450183c7650183c47501a206d98ec207e204c58fdd8e8216558e2338c14603c6950083c6850003c7a50083c7b5002206558e4207e2075d8f598e83c6d50003c7c50083c7e50083c4f500a206d98ec207e204c58fdd8e8216558e2334c14603c6150083c6050003c7250083c735002206558e4207e2075d8f598e83c6550003c7450083c7650083c57500a206d98ec207e205dd8dd58d8215d18d2330b146b14563e4bc006f20505f93841900058d630495016f20d05e13040a161395490022950c65aee8833d050093955400d29513965c00568597300000e78060f693954400a29513850a1613964c0097300000e78000f5231d3a21033501462330a13603358146833501470336814783dcaa212334a1362338b136233cc13613851c00b14563e4bc006f20704c33863b416304a6006f209057a66985098e04d2949385042213840a220e06228597300000e78020ef014593153500a2958c6133369501239ca5203295b3b6ac0093c61600758e23b8552165f2033581378335013703368136833601362334a1662330b166233cc1642338d1645285866763130b00568513060178ca85e2866a879770ffffe78080c7033501658335816503360166833681662330a15a2334b15a2338c15a233cd15a03350a21d687ee846e8cc66d6e8de31005d411a081494a6419e06f2090516a699770ffffe780c0c023380520231d052023308522930519002338a420231c04202ae92eed130da122930ba124630439016f20d04e8355a52129466374b6006f20904e1b861500231dc520139655008336015b2a960337015a8337815b14ea8336815a18e21cee1307052214e6139645002a96233096162334b6178505139635003a962330560123b8aa20239cba2039a8130601785285ca85e2866a879770ffffe78040b9130da122930ba124854d930a40088a7585052ef1327592757266d2662aeb2ee732e3b6fe280b0c1a1306200497300000e780a0d7034481177d461305111e9305911797300000e78040d6814c81491375e40f2300a11e05447e75de75233ca1203e751e762338b120667c2334a120a2e42330c120230031230949630a0c2a0a68e28283d8625b01451387825b93975800b30517013383f5001386725d63036706aa830345070293f5f90fb3b4a5002d8d3335a000b3059040c98d95e501541305f121b28421c88345050083c70400b3b6f500bd8db335b000b306d040d58dfd147d150504e5d1138513001307170213061602e385b5fb13f5f50f09cd631608003da4c683630508228e039e9283b282727d1885bf33855303169583458500930485006387052003c5b40183c5a40103c6c40183c6d40122054d8d4206e206558e518d83c5f40103c6e40183c6040203c71402a205d18dc2066207d98ed58d82154d8d233ca17803c5340183c5240103c6440183c6540122054d8d4206e206558e518d83c5740103c6640183c6840103c79401a205d18dc2066207d98ed58d82154d8d2338a17803c5b40083c5a40003c6c40083c6d40022054d8d4206e206558e518d83c5f40003c6e40083c6040103c71401a205d18dc2066207d98ed58d82154d8d2334a17803c5340083c5240003c6440083c6540022054d8d4206e206558e518d83c5740003c6640083c6840003c79400a205d18dc2066207d98ed58d82154d8d2330a17803c5b40383c5a40303c6c40383c6d40322054d8d4206e206558e518d83c5f40303c6e40383c6040403c71404a205d18dc2066207d98ed58d82154d8d2334a16603c5340383c5240303c6440383c6540322054d8d4206e206558e518d83c5740303c6640383c6840303c79403a205d18dc2066207d98ed58d82154d8d2330a16603c5b40283c5a40203c6c40283c6d40222054d8d4206e206558e518d83c5f40203c6e40283c6040303c71403a205d18dc2066207d98ed58d82154d8d233ca16403c5340283c5240203c6440283c6540222054d8d4206e206558e518d83c5740203c6640283c6840203c79402a205d18dc2066207d98ed58d82154d8d2338a16403c41400054931a8c9a403c4140093852400130501787d4697300000e78080a6014903c524046306052003c5d40583c5c40503c6e40583c6f40522054d8d4206e206558e518d83c5140603c6040683c6240603c73406a205d18dc2066207d98ed58d82154d8d233ca14603c5540583c5440503c6640583c6740522054d8d4206e206558e518d83c5940503c6840583c6a40503c7b405a205d18dc2066207d98ed58d82154d8d2338a14603c5d40483c5c40403c6e40483c6f40422054d8d4206e206558e518d83c5140503c6040583c6240503c73405a205d18dc2066207d98ed58d82154d8d2334a14603c5540483c5440403c6640483c6740422054d8d4206e206558e518d83c5940403c6840483c6a40403c7b404a205d18dc2066207d98ed58d82154d8d2330a14603c5d40783c5c40703c6e40783c6f40722054d8d4206e206558e518d83c5140803c6040883c6240803c73408a205d18dc2066207d98ed58d82154d8d233ca13603c5540783c5440703c6640783c6740722054d8d4206e206558e518d83c5940703c6840783c6a40703c7b407a205d18dc2066207d98ed58d82154d8d2338a13603c5d40683c5c40603c6e40683c6f40622054d8d4206e206558e518d83c5140703c6040783c6240703c73407a205d18dc2066207d98ed58d82154d8d2334a13603c5540683c5440603c6640683c6740622054d8d4206e206558e518d83c5940603c6840683c6a40603c7b406a205d18dc2066207d98ed58d82154d8d2330a13683ca3404054b29a883ca340493854404130501467d4697300000e7800084014b03358179833501790336817883360178233ca15a2338b15a2334c15a2330d15a033501658335816503360166833681662338a126233cb1262330c1282334d128033501468335814603360147833681472334a1222338b122233cc1222330d124033581378335013703368136833601362338a1762334b1762330c176233cd1740335815b8335015b0336815a8336015a233ca1782338b1782334c1782330d178033501278335812703360128833681282338a164233cb1642330c1662334d166033581228335012303368123833601242338a172233cb1722330c1742334d174033501778335817603360176833681752330a172233cb1702338c1702334d170139a8903cee893f9790009456312a9041355ba03ac1a2e9503450500335535010589930a4008630a052c1305015a7d46814597200000e780606388162c0b1306200497200000e780406f014a0149f1a1a28d230081469305017813060002130401781305114697200000e780006d9305016513060002930401651305114897200000e780806ba300614b2301514b93050173130600021305314a97200000e780c06993058170130600021305314c97200000e78080681355ba036e8aac1a2e95034505003355350105892c0b19e903498119034a91191304a1199304a11b9305114a03459401034684018346a4010347b4012205518dc2066207d98e558d0346d4018346c4010347e4018347f4012206558e4207e2075d8f598e0216518d233ca15a034514010346040183462401034734012205518dc2066207d98e558d034654018346440103476401834774012206558e4207e2075d8f598e0216518d2338a15a03459400034684008346a4000347b4002205518dc2066207d98e558d0346d4008346c4000347e4008347f4002206558e4207e2075d8f598e0216518d2334a15a034514000346040083462400034734002205518dc2066207d98e558d034654008346440003476400834774002206558e4207e2075d8f598e0216518d2330a15a03c5940003c6840083c6a40003c7b4002205518dc2066207d98e558d03c6d40083c6c40003c7e40083c7f4002206558e4207e2075d8f598e0216518d2330a17603c5140103c6040183c6240103c734012205518dc2066207d98e558d03c6540183c6440103c7640183c774012206558e4207e2075d8f598e0216518d2334a17603c5940103c6840183c6a40103c7b4012205518dc2066207d98e558d03c6d40183c6c40103c7e40183c7f4012206558e4207e2075d8f598e0216518d2338a17603c5140003c6040083c6240003c734002205518dc2066207d98e558d03c6540083c6440003c7640083c774002206558e4207e2075d8f598e0216518d233ca17488161306200497200000e780e044930a4008c669854d15a4034981199307a11903c5170083c5070003c6270083c6370022054d8d4206e206558e518d83c5570003c6470083c6670003c77700a205d18dc2066207d98ed58d82154d8d2330a15a03c5970083c5870003c6a70083c6b70022054d8d4206e206558e518d83c5d70003c6c70083c6e70003c7f700a205d18dc2066207d98ed58d82154d8d2334a15a03c5170183c5070103c6270183c6370122054d8d4206e206558e518d83c5570103c6470183c6670103c77701a205d18dc2066207d98ed58d82154d8d2338a15a03c5970183c5870103c6a70183c6b70122054d8d4206e206558e518d83c5d70103c6c70183c6e70103c7f701a205d18dc2066207d98ed58d82154d8d233ca15a9307a11b03c5970083c5870003c6a70083c6b70022054d8d4206e206558e518d83c5d70003c6c70083c6e70003c7f700a205d18dc2066207d98ed58d82154d8d2330a17603c5170183c5070103c6270183c6370122054d8d4206e206558e518d83c5570103c6470183c6670103c77701a205d18dc2066207d98ed58d82154d8d2334a17603c5970183c5870103c6a70183c6b70122054d8d4206e206558e518d83c5d70103c6c70183c6e70103c7f701a205d18dc2066207d98ed58d82154d8d2338a17603c5170083c5070003c6270083c6370022054d8d4206e20683c55700558e518d03c64700a20583c6670003c77700d18d034a9119c2066207d98ed58d82154d8d233ca174881613061002814597200000e7806015c66923042123a30441239305015a130600026a8597200000e780802093058175130600025e8597200000e780601f881c8c161306200497200000e780601e630c0920281d0c041306100297200000e780201d03451d0083450d0003462d0083463d0022054d8d4206e206558e518d83455d0003464d0083466d0003477d00a205d18dc2066207d98ed58d82154d8d2330a17803459d0083458d000346ad008346bd0022054d8d4206e206558e518d8345dd000346cd008346ed000347fd00a205d18dc2066207d98ed58d82154d8d2334a17803451d0183450d0103462d0183463d0122054d8d4206e206558e518d83455d0103464d0183466d0103477d01a205d18dc2066207d98ed58d82154d8d2338a17803459d0183458d010346ad018346bd0122054d8d4206e206558e518d8345dd010346cd018346ed010347fd01a205d18dc2066207d98ed58d82154d8d233ca17803c59b0083c58b0003c6ab0083c6bb0022054d8d4206e206558e518d83c5db0003c6cb0083c6eb0003c7fb00a205d18dc2066207d98ed58d82154d8d233ca16403c51b0183c50b0103c62b0183c63b0122054d8d4206e206558e518d83c55b0103c64b0183c66b0103c77b01a205d18dc2066207d98ed58d82154d8d2330a16603c59b0183c58b0103c6ab0183c6bb0122054d8d4206e206558e518d83c5db0103c6cb0183c6eb0103c7fb01a205d18dc2066207d98ed58d82154d8d2334a16603c51b0083c50b0003c62b0083c63b0022054d8d4206e206558e518d83c55b0003c64b0083c66b0003c77b00a205d18dc2066207d98ed58d82154d8d2338a164054b95a017a5feff93054552130600021305912297200000e780e03d8345012701254d8d05e117a5feff93052550130600021305112797200000e780c03b01256309055c281d0c041306100297200000e780e0f7130501787d46ea8597200000e780e0f6014be6e003450127630a05209307212703c5970183c5870103c6a70183c6b70122054d8d4206e206558e518d83c5d70103c6c70183c6e70103c7f701a205d18dc2066207d98ed58d82154d8d233ca14603c5170183c5070103c6270183c6370122054d8d4206e206558e518d83c5570103c6470183c6670103c77701a205d18dc2066207d98ed58d82154d8d2338a14603c5970083c5870003c6a70083c6b70022054d8d4206e206558e518d83c5d70003c6c70083c6e70003c7f700a205d18dc2066207d98ed58d82154d8d2334a14603c5170083c5070003c6270083c6370022054d8d4206e206558e518d83c5570003c6470083c6670003c77700a205d18dc2066207d98ed58d82154d8d2330a1469307212903c5970083c5870003c6a70083c6b70022054d8d4206e206558e518d83c5d70003c6c70083c6e70003c7f700a205d18dc2066207d98ed58d82154d8d2334a13603c5170183c5070103c6270183c6370122054d8d4206e206558e518d83c5570103c6470183c6670103c77701a205d18dc2066207d98ed58d82154d8d2338a13603c5970183c5870103c6a70183c6b70122054d8d4206e206558e518d83c5d70103c6c70183c6e70103c7f701a205d18dc2066207d98ed58d82154d8d233ca13603c5170083c5070003c6270083c6370022054d8d4206e206558e518d83c5570003c6470083c6670003c77700a205d18dc2066207d98ed58d8215034911274d8d2330a136854c29a803491127130501467d469305212797200000e780c0d3814c03358179833501790336817883360178233ca1342338b1342334c1342330d134033501658335816503360166833681662330a1322334b1322338c132233cd132033501468335814603360147833681472330a1302334b1302338c130233cd13003358137833501370336813683360136233ca12e2338b12e2334c12e2330d12e63030c028a642c1d62859770ffffe78000cd2e8471c5638604120e046294033c8472fd14cdb7900508622330a15608660c6a030686018334812b2334a1562338b156230cc1569770ffffe78040b2833501562a84233c955a033581562330b45c83350157233004002334a45c030581572338b45c8544231b945a230ca45c23046401a30444011305a4008c061306000297200000e78020c21305a4020c161306000297200000e78000c123059405a30524051305c4040c061306000297200000e78060bf1305c4068c151306000297200000e78040bea2fc02e1866c6f001002330554032a9c23046c01a3044c011305ac008c061306000297200000e780a0bb1305ac020c161306000297200000e78080ba23059c05a3052c051305cc040c061306000297200000e780e0b81305cc068c151306000297200000e780c0b7866c7daf4afc940588628c66906a83c686012330a1562334b1562338c156230cd156230cd1582338c1582334b1582330a15883596c5b0339812b2d4563f9a906da8dd28b13058c5b130b140093145400b3058500ae94330a540363fc69072380240113558903a383a400135509032383a40013558902a382a400135509022382a40013558901a381a400135509012381a40013558900a380a4001385840093050158654697200000e78000ad6da0930b4008054d914a154552f85af46369a4126303a412014d19456311a4120144954a39aa93155b005a952e9533848940131654002296a68597200000e780c0ed13558903a383a400135509032383a40013558902a382a400135509022382a40013558901a381a400135509012381a40013558900a380a400238024011385840093050158654697200000e78000a413058c00b305450133065b0332953306540397200000e78040e78529629a2304ba01a3047a011305aa008c061306000297200000e78080a01305aa020c161306000297200000e780609f23059a056275a305aa041305ca040c061306000297200000e780a09d1305ca068c151306000297200000e780809c231b3c5b854d6da463020c600a653384ad400c0462859770ffffe780209d630f05586305b45f8e05e29503bc85720504cdb7a28a19a06514994a9770ffffe780e0832a8b23300500231b055a83596c5b93c4faffce94231b955a930d8c5b93955a0033855d01aa95130501651306100297200000e7800095130a8c0033857a035295834b050093051500130501781306300897200000e780e092314563e4a4006f10a06c66f0ea8c138d1a003385a941630495006f10e07213058b5b93155d00ea9dee9513965400269697200000e780608f13064008b305cd02d29513058b003386c40297200000e780c08d231b5c5b1305015a930501651306100297200000e780408c13050146930501781306300897200000e780008b628d63930c005a8d83596d5b13058d5b930d140093145400b3058500ae94930a4008330a540363fab9052380240113558903a383a400135509032383a40013558902a382a400135509022382a40013558901a381a400135509012381a40013558900a380a4001385840093050158654697200000e780808359a093955d006e952e9533848940131654002296a68597200000e78080c613558903a383a400135509032383a40013558902a382a400135509022382a40013558901a381a400135509012381a40013558900a380a400238024011385840093050158654697100000e780c07c13058d00b305450133865d0332953306540397200000e78000c0854d027485296a9a22752304aa004275a304aa001305aa008c061306000297100000e780c0781305aa020c161306000297100000e780a07723058a046275a305aa041305ca040c061306000297100000e780e0751305ca068c151306000297100000e780c074231b3d5b130581759305015a1306100297100000e78040738816930501461306600897100000e7802072130da12209456397ab00930ba124866cc669b9a613058162930581751306100297100000e780a06f1305015a8c161306300897100000e780806e03350c00c669014a630705225a84835c4c5b2a8c13058170930581621306100297100000e780006c230071479305015a130630081305114697100000e780806a630400006f10804783596c5b2d4563eba92a52fc854d114a154522f8930b400863efac006389ac00814d19456397ac00814c154a29a0668a19a0e51c194a9760ffffe780e0532a8b23300500231b055a03596c5b9344faffca94231b955a930a8c5b93155a0033854a01aa95130581751306100297100000e780c06213048c0033057a032295034d05009305150088161306300897100000e780c060314563e4a4006f10803aee8b930d1a003305b941630495006f10603d13058b5b93955d00ee9ad69513965400269697100000e780605d930a4008b3855d03a29513058b003386540397100000e780c05b231b4c5b13050173930581751306100297100000e780405a130501788c161306300897100000e780205903546b5b13051400b1456364b4006f10c032338649416304a6006f104036627a050a8e0de29d93858d7293048b720e06268597100000e7808055014593153500a6958c6133368500239aa55a3295b336a40093c61600758e23b0650165f21305016e930501731306100297100000e780005213050165930501781306300897100000e780c0506285854dc66963930b005a851306817093060146e68542779760ffffe780c03e0945630fad10ea8b130581629305016e1306100297100000e780004d1305015a930501651306300897100000e780c04b03350c005a84e31e05dce67499e06f10e02d0a699760ffffe780c0372a8423300500231b055a233495721305190080e0239a045aa2fc2ae1130da122866c630449016f10402b8354645b2945637495006f10402b130984721b851400231ba45a13955400b30594002e951305855b930581621306100297100000e780e0433385540322952304750125059305015a1306300897100000e78020428504139534004a952330650123308b00231a9b5aa1a02300015a631eb40923308137233401362338b136130501468c161306015a9760ffffe780604759aa13068170930601466285e68522879760ffffe780e02cc669130da122866c930ba124aa64850426e57e75de753e769e762aeb2ee732e3b6fe280b90133414981cce8597a0ffffe78020af13f51c00631e0516a66413f5f40f130515f0933c1500138414008813ac1a26869750ffffe78080f0a6896fe0afe18e05e29503b5857219c8b30580400356655b0e06329503358572fd15edf98355655bfd152338a164233c01642330b16613050146930501651306015a9760ffffe780803b13050178930501461306500a97100000e780403103358150033a81518355655b03340151aa84636fba00046191c8035a455b83d5645b05042685e378bafe19a0228a2a8413155a00b38544012e959309855b33055a03269513098500881613061002ce8597100000e780c02b93050178130610024e8597100000e780a02a1306400813051138ca8597100000e7808029130640084a859305117a97100000e780602809cc0e0ad29483b404737d14c66919c483b484727d146dfc11a0c669130501468c161306500a97100000e780802523349150233801502a658345015a7d152ae5e38505e8667519e16f10200c8a6599e16f10400c03368572b2fcfd152ee12330060097f0feffe780a03285b5a8082c0b97a0ffffe78020b36fd00ff92689aa84033a8148833a014813155900229583459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18d233cb13683451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2338b13683459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2334b13683451500034605008346250003473500a205d18dc20662070346550083474500d98ed58d22065d8e834665000347750093174900b309f400c2066207d98e558e0216d18d2330b136930501781306000297100000e780000e03b5891683b5091623b0591723b4491791cc0e094a9403348422fd14930a400881c803340422fd14edfc19a0930a400803368137833601370337813683370136233cc1462338d1462334e1462330f1462330b1482334a14823388148233c01480a758345015a7d152af199e16fe0afad4a65e30d0570ea65e38f05700336052232e9fd152eed2338062097f0feffe780c0156fe04fabe6650676a6762eef467732f336f7e6753afb2a660a643339b000b3062041b3f9c600638d09063336200193361500758e11ca054909c483b585727d146dfc014a2e8521a02e8ae30a09668355655b6362b4020461e381045a0354455b050a97f0feffe780200f83d5645b2685e373b4fe26858145fd190504e3050afa0e042295033585729304faff81450144d9d803358572fd14edfc8145014461b7630a090219e52e8509c4033585727d146dfc0c6191c92e8497f0feffe780c0090c602285edf911a02a84228597f0feffe7808008ca6501450a766a6a3339b000b3062041b3f9c600638e09063336200193361500758e01ce054963070a0083b505227d1ae31d0afe81442e8521a0ae84e30c095a8355a5216363ba0203340521e306044e035a8521850497f0feffe780a0028355a4212285e372bafe22858145fd19050ad5d00e0a529503350522fd148145014ad1d803350522fd14edfc8145014a59b7630e090209e92e8563070a00033505227d1ae31d0afe8335052199c92e8497f0feffe78020fd833504212285e5f911a02a84228597f0feffe780c0fb13050004854597f0feffe78060fae3040558aa8dc26703c5970183c5870103c6a70183c6b70122054d8d4206e206558e518d83c5d70103c6c70183c6e70103c7f701a205d18dc2066207d98ed58d82154d8d233ca14603c5170183c5070103c6270183c6370122054d8d4206e206558e518d83c5570103c6470183c6670103c77701a205d18dc2066207d98ed58d82154d8d2338a14603c5970083c5870003c6a70083c6b70022054d8d4206e206558e518d83c5d70003c6c70083c6e70003c7f700a205d18dc2066207d98ed58d82154d8d2334a14603c5170083c5070003c6270083c6370022054d8d4206e206558e518d83c5570003c6470083c6670003c77700a205d18dc2066207d98ed58d82154d8d2330a146130501482c0b1306000297100000e78060d893050146130600046e8597100000e78040d785458546854c6e8501469770ffffe78080af6265033c050109452afa02fe82e2e3090c280949014b014482e46265033a05001795feff130565afaae893044006130d00108949b3058a0003c50500130685fba546e3eec62a0e06c66636961062930a14000286e36f2b23d27933059b024e950344e5fb130940068944e305943e1306c5f9835bc5f90355c6018355a6018356e6010357060242054d8d82164217d98e558d2334a1280355460183552601835666010357860142054d8d82164217d98e558d2330a1280355c6008355a60042058356e600035706014d8d9305360282164217d98e558d233ca126035546008356260003576600035686004205558d02174216598e518d2338a126130610041305117897100000e78080c523008178791bdae233052b034e95034425020949e3009434835405008355c5010356a5018356e50103570502c205d18d82164217d98ed58daee183554501035625018356650103578501c205d18d82164217d98ed58d2efd8355c5000356a500c2058356e500035705014d8e9305350282164217d98e558e32f9035645008356250003576500035585004206558e02174215598d518d2af5130610041305113697100000e78000bb33c574011335150093b50b106d8d23008136e307050ca8082c115e869740ffffe78020721305015a8c1c5e869740ffffe7802071a8089305015a1306000297100000e78020f90125e31c050813958b036d912c112e950345050093f57b003355b5000589630d056c13050146b008930601789816d9ad2665e314050626651a056e9583459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18d233cb14683451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2338b14683459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2334b14683451500034605008346250003473500a205d18dc2066207d98ed58d034655008346450003476500834775002206558e4207e2075d8f598e0216d18d2330b14683459503034685038346a5030347b503a205d18dc2066207d98ed58d0346d5038346c5030347e5038347f5032206558e4207e2075d8f598e0216d18d233cb13683451503034605038346250303473503a205d18dc2066207d98ed58d034655038346450303476503834775032206558e4207e2075d8f598e0216d18d2338b13683459502034685028346a5020347b502a205d18dc2066207d98ed58d0346d5028346c5020347e5028347f5022206558e4207e2075d8f598e0216d18d2334b13683451502034605028346250203473502a205d18dc2066207d98ed58d034655028346450203476502034575022206558e42076205598df276518d02154d8d2330a1366319db00081ada859790ffffe78080fe166bd27933059b023384a9002310040013052400930501461306000297100000e780808f23010402130534028c161306000297100000e780208e050bdae226650505aae4f9a133356001b3b58a016d8d630e055ed29a83ca0a0063940a00930a00107d1bdae233059b024e95834425026389247b835c05008355c5010356a5018356e50103570502c205d18d82164217d98ed58d233cb13683554501035625018356650103578501c205d18d82164217d98ed58d2338b1368355c5000356a500c2058356e500035705014d8e9305350282164217d98e558e2334c136035645008356250003576500035585004206558e02174215598d518d2330a136130501461306100497100000e780008103358137833501370336813683360136aaf8aef4b2f0b6ec2300917893050146130610041305117897000000e780007e63f7ac514675a6750676e666233ca15a2338b15a2334c15a2330d15a63820a2c8144b38b9c0013950b0341916371a54f1305015aac085e869740ffffe780603313958b036d91ac082e950345050093f57b003355b500058915c11305014613061002814597000000e780606a88161306015a93060146130701780da01305014613061002814597000000e780406888161306015a9306017813070146de859790ffffe78020e98504130501788c161306200497000000e7806072139504034191e36155f739ac63050b44930b140263e48b50636f7c43637d746133855b4193050002631eb55cb3055a01130600021305117897000000e780606e7d1bdae2d2792300017833059b024e958344250289456392b408cda3630d0b3e930b240463e18b4c63677c3f63f38a4d130524026360ac4c63e0ab5c130940063386ab4093060002631ed656d29a83c40a0013842500b305aa00130600021305217a97000000e780c0671306000213052178a28597000000e780a0667d1bdae2d279a30091782300917933052b034e958344250289456388b456035405008355c5010356a5018356e50103570502c205d18d82164217d98ed58daef883554501035625018356650103578501c205d18d82164217d98ed58daef48355c5000356a500c2058356e500035705014d8e9305350282164217d98e558eb2f0035645008356250003576500035585004206558e02174215598d518daaec130610041305113697000000e780c05b230091366374a42f1305015aac0822869740ffffe780a013131584036d91ac082e9503450500937574003355b500058909c9130501461306015a93060178981601a8130501461306015a941613070178a2859790ffffe780a0cb930440067275631cab000949081ada859790ffffe78060c1166bd27911a00949050433059b02b384a90023908400138524009305015a1306000297000000e78000521385240293044006930501461306200497000000e7808050050bdae2de8ae5a8e68b0335015a8335815a0336015b8336815b2330a1362334b1362338c136233cd13613050146930501781306200497000000e780a04c7275631aab00081ada859790ffffe78040b8166bd279854c93044006930a2400850b33059b023384a90023107401130524008c161306000297000000e780a04813052402930501461306200497000000e7806047166b9da013050146b008941613070178de859790ffffe78040bb930440067275631aab00081ada859790ffffe78020b1166bd279850b33059b023384a9002310740113052400ac081306000297000000e780204213052402930501461306200497000000e780e040050bdae2568463ed8aed05456319ab1252740355040013450510a66593c515004d8d631e051093052402130511659790ffffe780c0cf727511c5228597e0feffe780804d6e8597e0feffe780e04c03156165831541650356216583061165231aa172c205d18d033581662328b1728305016703348165233ca174833401662300b1762304d1221305912293050173194697000000e780603713558403230ba12213550403a30aa12213558402230aa12213550402a309a122135584012309a12213550401a308a122135584002308a122a307812213d58403230fa12213d50403a30ea12213d58402230ea12213d50402a30da12213d58401230da12213d50401a30ca12213d58400230ca122a30b91221305f12393058175254697000000e780c02e281413060002a26597000000e7804070814c01251334150005a0854c727511c5527597e0feffe780003d6e8597e0feffe780603c13044002e265886511c5886197e0feffe780203b6685a2850d618330817e0334017e8334817d0339017d8339817c033a017c833a817b033b017b833b817a033c017a833c8179033d0179833d81781301017f8280a308a16441bfad452685ada0b1459da097e0feffe780a0351785feff1305257c09a897e0feffe78080341785feff1305057b9305b00291a81795feff130595929305500399a01795feff1305358f25a81795feff1305958e3da01785feff1305e57a29a01785feff1305457af14531a85685e2859730ffffe780e00200001795feff1305b58b930580029720ffffe780207800001785feff1305657459bf1795feff1305a58493050003c5b71785feff1305e56e93050002c9bfad4566855dbf1795feff130595877dbf1795feff1305f58655bf1785feff1305657099bf1785feff1305c56fb1b71785feff1305256f89b71795feff130565829305100271b7ad454e8585bf1795feff13053583a5bf1785feff1305a56c29bf1785feff1305e57fe1bf1785feff1305656b19b71785feff1305a57b85bf1785feff1305256695bf13050002930500022db797e0feffe780602300001785feff13054568d1bd1785feff1305a567e9b51785feff13050567c1b55685de85f5bd1785feff1305056645bd1785feff130565655db571c693f7f50f2300f5003307c500a30ff7fe894663fcc60aa300f5002301f500230ff7fea30ef7fe994663f1c60aa301f500230ef7fea14663fac60893f5f50f9b9785003307a0400d8bad9f198e9b950701ad9f2a97719a1cc3b305c70023aef5fe63f5c6065cc31cc723aaf5fe23acf5fee14663fcc604137847005cc71ccb5ccb1ccf6108939807029396070293d8080223a2f5fe23a4f5fe23a6f5fe23a8f5fe33060641fd474297c69663f0c7020116937706fe93870702ba9714e314e714eb14ef13070702e31af7fe8280397122fc26f84af44ef052ec56e85ae45ee093f735006387074069c2aa8719a06303062a83c60500850513f735002380d7007d1685076df793f637003e87cdea3d48637dc804930806ff6378180133e8b700137878006304083093d84800138f1800120f2e9f2e87be86832e0700032e4700032387000328c70023a0d60123a2c60123a4660023a606014107c106e31eeffc85089208c695c6973d8a137886001377460093762600058a630c080083a8050003a84500a107a10523ac17ff23ae07ff11c798419107910523aee7fe6391061e09c603c705002380e7006274c27422798279626ac26a226b826b216182807d476379c70a094883c805009841638806290d486386061d9306c6fe03c3150003c8250093f306ff13843700938435009382330123801701a38067002381070113d94600ae92a687a28803a8170083a5570083a697001b53870103a7d7009b1f88001b9f85009b9e86001b5888019bd585019bd686011b1e87003363f3013368e801b3e5d501b3e6c60123a0680023a2080123a4b80023a6d800c107c108e39657fa9307190092073516b385f40033067640a29793780601137886009376460013772600058a6384080883cb050003cb150083ca250003ca350083c9450003c9550083c4650003c4750083c3850083c2950083cfa50003cfb50083cec50003ced50003c3e50083c8f50023807701a380670123815701a381470123823701a382270123839700a383870023847700a38457002385f701a385e7012386d701a386c70123876700a3871701c105c1076304080483c2050083cf150003cf250083ce350003ce450003c3550083c8650003c8750023805700a380f7012381e701a381d7012382c701a382670023831701a3830701a105a1079dc203c3050083c8150003c8250083c6350023806700a380170123810701a381d70091059107e30307e283c6050003c715008907238fd7fea38fe7fe890539b513f73700e31d07ec39b59306c6fe93f306ff1384170093841500938213012380170113d94600ae92a687a28803a8370083a5770083a6b7001b53870003a7f7009b1f88011b9f85019b9e86011b5888009bd585009bd686001b1e87013363f3013368e801b3e5d501b3e6c60123a0680023a2080123a4b80023a6d800c107c108e39657fa9307190092073d16b385f40033067640a297a1b593d84800938e18002e88033e88000333080085062334c7012330670041084107e3e5d6ff85089208c695c6973d8a01bb9306c6fe03c8150093f306ff13842700938425009382230123801701a380070113d94600ae92a687a28803a8270083a5670083a6a7001b53070103a7e7009b1f08011b9f05019b9e06011b5808019bd505019bd606011b1e07013363f3013368e801b3e5d501b3e6c60123a0680023a2080123a4b80023a6d800c107c108e39657fa9307190092073916b385f40033067640a29749b3aa8709b919ca0347050083c705007d166317f700050585057df6014582800345050083c705001d9d8280aa862e87b287630db50cb388c5403308c040b388a84006082e832a8e6372181b3346b5001d8a637fb50a63010612cdcb1386f7ff9d4563f8c51813061700b305c54093b5750093c5150093f5f50f638a0516b365e5009d896395051693f587ffba95033603002103210e233ccefee39a65fe13f687ff13f57700aa87b385c600329739cd0345070005462380a5006389c704034517000946a380a5006382c704034527000d462381a500638bc702034537001146a381a5006384c7020345470015462382a500638dc700034557001946a382a5006386c700834767002383f5003685828029ea3306f5001d8a65ca1386f7fffdd7b307c5007d5821a07d16e30106ffb305c70003c5050093f57700fd17a380a700e5f59d4763fac70ab2871d48e117b305f7008861b385f60088e1e369f8fe93777600cdd7fd173306f700834506003386f6002300b600f5b71376750041ca9385f7ffc9d72a867d5821a0fd15e38005f903450700050693777600a30fa6fe0507edf79d4763fcb704938885ff93f888ffa10833051601ba8703b807002106a107233c06ffe31aa6fe469793f77500130617008ddfba9711a005060347f6ff0505a30fe5fee31af6fe36858280cdba3685d5b713061700f9bfb287a5b73285ae8713061700e1f919b73e8625bf2a86be8549bfcdccccccccccccccd182e6ad7f520e5108c9bcf367e6096a1f6c3e2b8c68059b3ba7ca8485ae67bb6bbd41fbabd9831f2bf894fe72f36e3c79217e1319cde05bf1361d5f3af54fa54b598638d6c56d340101010101010101ff00ff00ff00ff00fffefefefefefefe80808080808080800a0a0a0a0a0a0a0aaf47e17a14ae4701555555555555555533333333333333330f0f0f0f0f0f0f0f01010101010101019a999999999999010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000088ab0a000000000000100000000000000400000000000000889b020000000000001008000000000040000000000000000100000000000000c0090100000000000000000000000000011101250e1305030e10171b0eb44219110112060000023901030e0000032e001101120640186e0e030e3a0b3b053f198701190000041101250e1305030e10171b0eb44219110155170000052e006e0e030e3a0b3b05200b0000062e001101120640186e0e030e3a0b3b050000072e006e0e030e3a0b3b0b200b0000082e011101120640186e0e030e3a0b3b0b360b0000091d00311311011206580b590b570b00000a1d0031135517580b590b570b00000b1d00311311011206580b5905570b00000c1d0031135517580b5905570b00000d2e006e0e030e3a0b3b0b3f19200b00000e2e011101120640186e0e030e3a0b3b0b3f1900000f1d0131135517580b590b570b0000101d01311311011206580b590b570b0000111d01311311011206580b5905570b0000121d0131135517580b5905570b0000132e006e0e030e3a0b3b053f19200b0000142e011101120640186e0e030e3a0b3b05360b3f190000152e011101120640186e0e030e3a0b3b053f190000162e0111011206401831130000172e0011011206401831130000182e001101120640186e0e030e3a0b3b0b0000192e011101120640186e0e030e3a0b3b0b00001a2e011101120640186e0e030e3a0b3b0500001b2e001101120640186e0e030e3a0b3b0b3f1987011900001c2e006e0e030e3a0b3b0b870119200b00001d2e011101120640186e0e030e3a0b3b05360b3f198701190000004d00000004000000000008019c2b00001c0023460000000000005213000024650100000000000e000000029b2f000002000000000324650100000000000e0000000152494f000050380000010b020000002326000004000000000008049c2b00001c00811700005c0000005213000000000000000000007011000002621a00000284050000052f0d0000b717000002f9050106aea2010000000000020000000152c8350000dd0c000002eb0102813f0000028333000005d23800003f2500000693030105d23800003f2500000693030105d23800003f2500000693030105d23800003f2500000693030105d23800003f2500000693030105cb2a0000932300000693030105122d0000944900000693030105a63b00005b3a00000693030105770c0000f90300000636050105d23800003f250000069303010000025f0d0000028333000005844200003f2500000801040105844200003f2500000801040105844200003f2500000801040105844200003f2500000801040105844200003f25000008010401059c330000b41800000801040105ff0b0000c137000008010401000005a60000003c4a00000273040105241400002d4400000273040105e7480000900500000249050105b8080000cc00000002490501053c2a0000f90300000261060100027f3300000282130000027c34000007ca4b00007b29000003d001000251410000075d1400008b490000038e01077b3e00007f330000038901077b3e00007f330000038901000002214c0000027631000008b0a2010000000000420100000152231700006238000005d303096500000020a30100000000000200000005f1360a161c00000000000005f115097200000032a30100000000000200000005f2360a231c00004000000005f215097f0000007aa30100000000000200000005fd360a301c00007000000005fd1509f300000088a30100000000000200000005fd470b00010000a2a3010000000000020000000503011e0b8c000000b4a301000000000002000000050701360c3d1c0000a0000000050701150b0d010000c2a301000000000002000000050701470b1a010000d0a301000000000006000000050f0133000002550c0000076e2d0000ac3e0000054301076b1b0000f204000005430107e8160000db10000005430107d1300000752b00000543010002512b00000d281500007f1d000005870100024e4700000d884a0000093c0000052a0100029d1500000e70ab010000000000700000000152163100007f330000059a0fd902000020090000059b11108c1d000076ab01000000000008000000054e1d11f71c000076ab010000000000080000001af80209094101000076ab010000000000080000001cef5000000a0f0300005009000005511c093c22000088ab01000000000004000000055116092103000096ab010000000000080000000551280fd724000080090000056514125b1e0000b0090000225901090a481e0000e0090000181209000000000002c60700000d5f3500007f1d000005870100020f0f00000e48b20100000000007200000001521c2900007f330000059a0fe5020000100e0000059b1110e01d00004eb201000000000008000000054e1d11f71c00004eb2010000000000080000001af8020909410100004eb2010000000000080000001cef5000000afa030000400e000005511c094922000064b20100000000000400000005511609b11b000070b201000000000008000000054f190fe4240000700e000005651412671e0000a00e0000225901090a481e0000d00e00001812090000000000020e4800000ebab2010000000000720000000152724800007f330000059a0ff1020000000f0000059b1110ed1d0000c0b201000000000008000000054e1d11f71c0000c0b2010000000000080000001af802090941010000c0b2010000000000080000001cef5000000a0f030000300f000005511c0956220000d6b20100000000000400000005511609b11b0000e2b201000000000008000000054f190ff1240000600f000005651412731e0000900f0000225901090a481e0000c00f0000181209000000000002210800000ee4b30100000000007000000001521f0300007f330000059a0ffd02000080100000059b1110fa1d0000eab301000000000008000000054e1d11f71c0000eab3010000000000080000001af802090941010000eab3010000000000080000001cef5000000afa030000b010000005511c0963220000fcb30100000000000400000005511609210300000ab4010000000000080000000551280ffe240000e0100000056514127f1e000010110000225901090a481e00004011000018120900000000000002a44d000013e90a00001e0b000009bd0601137f0300007a31000009f6060113964c00001944000009100701056b0d000088050000096e050114f2a3010000000000e4010000015289020000b834000009de04030b6206000010a40100000000000c00000009e504130b6f0600002ca40100000000000400000009ea04190b7c06000068a401000000000002000000090a051a1289060000d000000009170524112f20000050a50100000000000400000009800512111c20000050a5010000000000040000000fc702090b8222000050a5010000000000020000000f6d020c000000121b13000010010000091a0511123c2000004001000009940412121c200000700100000fc702090c82220000a00100000f6d020c0000001218220000d0010000090b05200b50010000e2a401000000000006000000149403160b6a010000f6a4010000000000040000001495030900122522000000020000090c05210b5d010000e8a401000000000004000000149403160b77010000faa4010000000000040000001495030900118906000014a50100000000001a000000090e0524112f2000001aa50100000000000400000009800512111c2000001aa5010000000000040000000fc702090b822200001aa5010000000000040000000f6d020c00000011d42000003ea40100000000001c00000009eb0416106f2000003ea40100000000001c00000013310910632000003ea40100000000001c00000012200910c71f00003ea40100000000001c00000012874c103a1f00003ea40100000000001c000000115331116d1f00003ea40100000000001c0000000b940d09109d1f00003ea40100000000001c0000000d3211102d1f00003ea40100000000001c000000107c09125a1c0000300200000bb0091d109c1c00004aa4010000000000020000000a2b3509270100004aa4010000000000020000000a5352000012af1f0000800200000bb1091510dd1f00004ca40100000000000800000010541c10802000004ca401000000000008000000115016092b2100004ca40100000000000800000012871f0000097e1f000056a40100000000000200000010541500000000000000000000152ca6010000000000780300000152454b00000c310000093c0512f6220000b0020000093e05170ce9220000e00200001583020f0011862100005aa6010000000000040000000947052511792100005aa60100000000000400000017410333110a1d00005aa6010000000000040000001708032711a81c00005aa6010000000000040000001ae5020909990000005aa6010000000000040000001c62500000000011541f00005ea6010000000000da0000000947052311471f00005ea60100000000006e0000000b8b010912f2200000100300000b5801100fe020000040030000138c190f3721000070030000132c12095a1c000082a6010000000000040000000c260e094f2100009aa6010000000000040000000c3212095b210000a6a60100000000000a0000000c39130967210000bca60100000000000a0000000c4125094321000096a6010000000000040000000c2e1000000011492000007ea6010000000000040000000b570112111c2000007ea6010000000000040000000fc702090b822200007ea6010000000000020000000f6d020c00000011f2200000eaa60100000000004e0000000b8c010910e0200000eaa60100000000004a000000138c191037210000eaa60100000000004a000000132c12095a1c0000eaa6010000000000040000000c260e096721000022a70100000000000c0000000c4125095b21000016a7010000000000040000000c3913094f21000012a7010000000000040000000c321200000000129f210000a0030000094c051312c4210000d003000017b90109119321000038a7010000000000120000001914010c10171d00003ea70100000000000400000017dc1f0b121e00003ea7010000000000040000001a5a010f000000000c0323000000040000094c051c11d42000006ca70100000000007201000009590523106f2000006ca701000000000072010000133109106320000072a70100000000001e00000012200910c71f000072a70100000000001e00000012874c103a1f000072a70100000000001e000000115331116d1f000072a70100000000001e0000000b940d09109d1f000072a70100000000001e0000000d3211102d1f000072a70100000000001e000000107c09125a1c0000300400000bb0091d109c1c00007ea7010000000000020000000a2b3509270100007ea7010000000000020000000a5352000012af1f0000800400000bb1091510dd1f000080a70100000000000800000010541c108020000080a701000000000008000000115016092b21000080a70100000000000800000012871f0000097e1f00008aa70100000000000200000010541500000000000000108d20000090a70100000000004e01000012220910241d000090a701000000000014000000123a270b8401000090a7010000000000060000001ad60d1f113e1d000096a7010000000000080000001ada0d200b311d000096a7010000000000080000001a460617000b4b1d00009ea7010000000000060000001adb0d24001063200000a4a70100000000001a00000012471510c71f0000a4a70100000000001a00000012874c103a1f0000a4a70100000000001a000000115331116d1f0000a4a70100000000001a0000000b940d09109d1f0000a4a70100000000001a0000000d3211102d1f0000a4a70100000000001a000000107c09125a1c0000b00400000bb0091d109c1c0000aea7010000000000020000000a2b350927010000aea7010000000000020000000a5352000012af1f0000000500000bb1091510dd1f0000b0a70100000000000800000010541c1080200000b0a701000000000008000000115016092b210000b0a70100000000000800000012871f0000097e1f0000baa701000000000002000000105415000000000000001063200000c0a70100000000001c00000012473510c71f0000c0a70100000000001c00000012874c103a1f0000c0a70100000000001c000000115331116d1f0000c0a70100000000001c0000000b940d09109d1f0000c0a70100000000001c0000000d3211102d1f0000c0a70100000000001c000000107c09125a1c0000300500000bb0091d109c1c0000cca7010000000000020000000a2b350927010000cca7010000000000020000000a5352000012af1f0000800500000bb1091510dd1f0000cea70100000000000800000010541c1080200000cea701000000000008000000115016092b210000cea70100000000000800000012871f0000097e1f0000d8a70100000000000200000010541500000000000000109920000012a801000000000012000000125a12096f2300001ea801000000000004000000127f0e0010e51c000040a80100000000000600000012501910651d000040a8010000000000060000001c1a0e11b41c000040a8010000000000060000001ae5020909a600000040a8010000000000060000001c62500000000a661c0000b00500001250190aa5200000f005000012541b0f721c00006006000012631a10c01c0000b2a8010000000000020000000a2b350934010000b2a8010000000000020000000a5352000009b1200000b4a80100000000000c00000012641b10bd200000caa801000000000012000000126616097c230000d6a801000000000004000000127f0e0009581d00003ca801000000000004000000124f2c10d21c000028a801000000000010000000124a1211d122000034a8010000000000040000001ccb051b11c322000034a8010000000000040000000e7e04080bb122000034a8010000000000040000000e2e03090000000000001289060000b006000009630528112f2000003aa90100000000000400000009800512111c2000003aa9010000000000040000000fc702090b822200003aa9010000000000020000000f6d020c000000111b13000066a90100000000002600000009650515123c200000f006000009940412121c200000200700000fc702090c82220000500700000f6d020c000000000d773b00002b30000009f20113bf180000642d000009f4050113fe330000442b00000943070105e8280000111e0000099c040116a2b10100000000009800000001520813000011ca190000aeb10100000000001800000009e6071b0b0b120000aeb10100000000000c0000001f170112001167180000d4b10100000000005800000009e8070911ab240000deb10100000000004a0000001f650127115b170000e0b10100000000004800000020270516116f170000f4b1010000000000060000001f66013c0b6f060000f4b1010000000000060000001f700109000b0b120000fcb1010000000000140000001f6701150b0b12000012b2010000000000160000001f6901110000000013db0700002525000009e507010002ec1b000005801800000e3200000993040100021432000002b834000006d6a5010000000000560000000152544d0000a61b000009f304000005ac090000104d000009640401053e100000d10900000979040115b2a90100000000007e0100000152803c00000e3200000938040cff110000800700000939041912f71f0000b0070000094d041d0a7e1c0000e00700001d2f1100124f130000100800000956041a115c1300003aaa01000000000018000000096b04150bb301000040aa010000000000120000000981042c00115c13000060aa01000000000018000000096c04190bb301000066aa010000000000120000000981042c0011721d000080aa010000000000040000000973041f111e1e000080aa010000000000040000001a96011a09b300000080aa0100000000000400000018ee1c00000bbf01000084aa010000000000080000000976040b00120320000040080000093f041d0a8a1c0000700800001d2f11000bcb010000d2aa0100000000000a00000009460415127f1d0000a0080000095d0426122a1e0000e00800001a5a010f10361e000000ab0100000000000400000018d93609c000000000ab0100000000000400000018ee1c0000000002f101000007fa3f0000f83b00001f550102273b00000ee0ab010000000000bc01000001526a380000642d00001f1f0f17210000100a00001f20121204210000400a0000133f0509110322000066ac010000000000d40000001372020f11a61d000070ac01000000000008000000249e01320b911e000070ac010000000000080000001a5a01090011db1e000078ac010000000000ac00000024a2012209e71e00007eac0100000000001a000000252c1010f31e000098ac0100000000008c000000252f0510cd00000098ac0100000000000c0000002552160b8401000098ac0100000000000c0000000640051600100b1f0000deac0100000000000a000000256a160996230000deac010000000000020000002514070010ff1e0000c8ac0100000000000a0000002569160989230000c8ac010000000000020000002514070009da000000bcac0100000000000400000025651b09e71e000010ad0100000000001400000025771609e71e0000f0ac01000000000012000000255a1e000011b31d000030ad0100000000000200000024b701430b911e000030ad010000000000020000001a5a01090011a222000032ad0100000000000400000024b8011c11c81e000032ad010000000000040000000ea9050d09aa1e000032ad01000000000004000000231a0900000000000fac210000700a00001f252712f0210000a00a0000175f040d12dd210000d00a00002445022912991d0000000b000024de0309119522000042ac0100000000000a0000001a09091311bc1e000042ac0100000000000a0000000ea9050d09aa1e000042ac0100000000000a000000231a0900000000000000000287400000020848000005920400007b2900001f3501010002641b000005ca2400007b2900001f6501010000026a2b000005144d0000294a00001f6f01011582af0100000000002001000001526f0a0000084800001f34011291240000b00b00001f3501231148170000a6af010000000000de00000020270516126f170000e00b00001f3601100c6f060000100c00001f700109000b0b120000ceaf010000000000160000001f3801150c0b120000400c00001f4101110bbe24000004b0010000000000020000001f410111127a180000700c00001f3c01220f25120000b00c00001f1a09119118000024b00100000000000a00000009a30412091023000024b00100000000000a0000001f1a260000000b0b12000070b0010000000000120000001f3e0111000000138b1e0000641b00001f6301010002304b000007501e0000363000001f15010002a3090000023630000007f73700007b2900001f1a01000002591b0000053b300000ec0400001f7b010105cf0e0000294a00001f9101010002de4c000002ec04000005773000007b2900001f7c0101000002c83a000015a2b00100000000000001000001524b050000ec0400001fd40112a4180000f00c00001fd50109129e240000200d00001f7c012311c9180000deb0010000000000c40000002027051612b1180000500d00001f7d01100c6f060000800d00001f920109000b0b120000f2b0010000000000180000001f8801150b0b12000018b1010000000000180000001f7f0115127a180000b00d00001f8301220f25120000e00d00001f1a09119118000044b10100000000000a00000009a30412091023000044b10100000000000a0000001f1a260000000b0b1200008cb1010000000000160000001f85011100000000000541340000ba2400001f1301010002fb320000169cad010000000000b400000001523c1a00001015260000aaad0100000000009600000009a41a1103260000aaad010000000000960000002679022a0cf6250000300b000026b6060f0000001750ae010000000000380000000152481a000007d51900000133000009a30107d74700001e4f000009bf010002833300001888ae0100000000000a0000000152744b00003a45000009c61992ae010000000000b60000000152654500000133000009ca103c1a0000a0ae010000000000a200000009cb091015260000a2ae0100000000009600000009a41a1103260000a2ae010000000000960000002679022a0cf6250000700b000026b6060f000000001948af0100000000003a0000000152d13a00001e4f000009ce09481a000068af0100000000001400000009cf090000022a0a000005011100007f33000009bb09010002d30c00001a2cb3010000000000160000000152373300004c11000009d0080b0e1b00002cb30100000000001600000009d0083e00000002c73c0000029b4d0000021a4c0000199ca2010000000000040000000152340a0000824f000001fa10a10100009ca20100000000000400000001fa0509340000009ca20100000000000200000003d21e00000000024b2f000002d007000005512f0000d71000002742020100000002872900001ba0a20100000000000e0000000152190f00003b4b000004341ba4a90100000000000e00000001525417000010310000046e1c36400000301300000495011c68100000373400000485010002cb3c000005ab0a0000b5110000075f0a0105ab0a0000b5110000075f0a0105ab0a0000b5110000075f0a0105ab0a0000b5110000075f0a0100028934000002c81e000002472500000752360000d14800000a7c0107013e0000c10100000a7c0107982c00004c4400000a7c0107384e0000304100000a7c0107c71c0000dc3f00000a7c010002243900000712000000cb1b00000a4b0107a82f0000d64c00001c5b0107cd340000a32300001c5b0107b3230000373700000a4b0100022e4e000005db3900004c4400001cc7050100028333000007740b0000eb3d00001c190100024d0c000007411d0000024500001cd9010000028333000005b1120000f81b00001ae4020105771c00002d2a00001a56010105034700005d4a00001acb0d010553270000d14000001a9806010518060000e84000001a4206010568440000620900001a860d01056b2a0000b72a00001a16040105303b0000da3d00001ae4020105db1a0000f81200001a8f010105bc440000563200001a56010105ed270000da0900001af70201055b0e0000521900001a040901054c040000311b00001a560101054c040000311b00001a56010102b6070000033ab20100000000000e0000000152bd450000b53c00001a0b0d0005ed270000da0900001af7020105ed270000da0900001af7020105ed270000da0900001af702010002b403000002273b000007af050000c534000018d701074d3700001d2b000018e30107f20d00002613000018d701075a410000ea33000018e3010002653a000005fa010000b149000018ec01010002833300000767320000f41800001811010767320000f41800001811010767320000f41800001811010767320000f41800001811010002874000000510160000c5340000185f01010000029e0d000002de4c000007a7150000d33e000023520100028333000007851d00007c40000023190107851d00007c4000002319010000022f30000007601900002f30000025290107e13e0000193f00002534010def4a0000021e00002547010799100000ce4100002513010799100000ce410000251301000002c81e000002a12f000002dd2b0000025b4600000585130000522500000baa0901058b3f0000d24200000b8f0d010567390000f60000000b56010105ec080000dd0f00000b8a0101000002cd11000002d31100000791290000d63c00000d310102670d000007a5430000dd1100000d35010000000002334a0000028431000002273b00000788310000cd1e00001078010002b54d00000770460000ea200000105401000002ae4d000002273b0000072b080000c5130000114d01020c00000002da48000007cc170000590000001150010000000002bd1c000002a30900000763060000a92700001d2e010793140000fa2300001d2e0100000002df08000002273b0000050e490000982200000f6c02010002474a000005a92200004c4400000fc6020105a92200004c4400000fc6020105a92200004c4400000fc602010000000208000000020c0000000d280b0000b31b0000128601074a0f000064460000121a0102b31b0000078c2000007b290000128701000d2b090000cc1a000012260107f54000004a140000127a0107512c0000d201000012720107512c0000d201000012720107f54000004a140000127a010002c81e0000028333000007254c00000c00000013300107be4d00001f0100001329010002de4c000007011c00001f010000138a010002e2320000053e280000620c0000136c0201000230450000050f2e0000f0320000133e0501000002680b00000790400000ca3f00000c180107e62b0000ae3900000c240107ff0f0000252c00000c0b01073e230000802300000c1101073e230000802300000c1101073e230000802300000c11010002833300000529390000cf3600001707030105e7290000504a00001740030107a80d0000352c000017d30105d53600001137000017b80101050a0400006c400000175b04010002a12f000002933300000524010000ab05000019130101000002da4a000002512b000005b24e0000e24a000024dd03010002474a0000058c280000e24a00002441020100028333000005912e000012350000249b010100000002e348000005a23d0000de1b0000148f0301058f3400007e0f0000148f030102a92d0000029115000005804700007e4a000021e8010105804700007e4a000021e8010105804700007e4a000021e8010105804700007e4a000021e80101000000029e0d000002a20d000002ec00000005671a0000cc3600000e5305010002b1240000050f3c00005b2b00000ea80501050f3c00005b2b00000ea80501000005584700001d3200000e93040102573a000005e74c0000462c00000e2a030100057e090000462c00000e7d04010002e5080000028c33000005a00f00009c0500001556020105c6460000cb3d00001582020105ba0300005844000015bb030105f6060000a70e000015120601001d62ab0100000000000e000000015251420000a73c0000158b070311041c000064ab0100000000000c000000158c070509f81b000064ab0100000000000c00000004860500000002214c0000024e47000005e32f0000714a00001be4040105e32f0000714a00001be4040105e1490000114f00001bcd040105e1490000114f00001bcd04010000022c1b000002e32700001530ab010000000000120000000152184800007f3300001ebb02111812000030ab010000000000120000001ebc021b11dd14000030ab0100000000001200000009440709090b12000030ab010000000000120000001f59120000000002083500001542ab010000000000120000000152c20200007f3300001ed602111812000042ab010000000000120000001ed7021b11dd14000042ab0100000000001200000009440709090b12000042ab010000000000120000001f5912000000000002211500000354ab0100000000000e0000000152180500004413000020720602294b0000051d350000081a00002025050105320700006e3a0000202505010574070000263f00002025050100022d33000005e14100000d0a0000209b07010000023828000002481900000531240000b62d0000225801010531240000b62d0000225801010531240000b62d0000225801010531240000b62d00002258010100022d3300000e42b3010000000000a20000000152541100007f33000022830f08130000f00f000022830a12ca1900002010000009e6071b0c0b120000501000001f17011200116718000080b30100000000005800000009e8070911ab2400008ab30100000000004a0000001f650127115b1700008cb30100000000004800000020270516116f170000a0b3010000000000060000001f66013c0b6f060000a0b3010000000000060000001f700109000b0b120000a8b3010000000000140000001f6701150b0b120000beb3010000000000160000001f6901110000000000000002f106000002ef37000005082f00009119000026990601059a1900003b2f000026b5060102833300000599160000cb4700002677020100000000002c0000000200000000000800ffffffff24650100000000000e0000000000000000000000000000000000000000000000ec0100000200510000000800ffffffff9ca20100000000000400000000000000a0a20100000000000e00000000000000aea20100000000000200000000000000b0a20100000000004201000000000000f2a3010000000000e401000000000000d6a501000000000056000000000000002ca60100000000007803000000000000a4a90100000000000e00000000000000b2a90100000000007e0100000000000030ab010000000000120000000000000042ab010000000000120000000000000054ab0100000000000e0000000000000062ab0100000000000e0000000000000070ab0100000000007000000000000000e0ab010000000000bc010000000000009cad010000000000b40000000000000050ae010000000000380000000000000088ae0100000000000a0000000000000092ae010000000000b60000000000000048af0100000000003a0000000000000082af0100000000002001000000000000a2b00100000000000001000000000000a2b101000000000098000000000000003ab20100000000000e0000000000000048b20100000000007200000000000000bab201000000000072000000000000002cb3010000000000160000000000000042b3010000000000a200000000000000e4b301000000000070000000000000000000000000000000000000000000000022a301000000000026a30100000000002aa301000000000032a30100000000003ea301000000000042a30100000000000000000000000000000000000000000034a30100000000003ca301000000000042a30100000000004aa3010000000000000000000000000000000000000000007ca301000000000088a30100000000008aa301000000000094a301000000000000000000000000000000000000000000b6a3010000000000c2a3010000000000c4a3010000000000cca3010000000000000000000000000000000000000000006ca401000000000072a401000000000076a40100000000007ca401000000000030a501000000000060a50100000000000000000000000000000000000000000090a5010000000000b0a5010000000000d0a5010000000000d6a50100000000000000000000000000000000000000000098a5010000000000a0a5010000000000d0a5010000000000d6a50100000000000000000000000000000000000000000098a5010000000000a0a5010000000000d0a5010000000000d6a50100000000000000000000000000000000000000000098a5010000000000a0a5010000000000d0a5010000000000d6a501000000000000000000000000000000000000000000e2a4010000000000e8a4010000000000f6a4010000000000faa401000000000000000000000000000000000000000000e8a4010000000000eca4010000000000faa4010000000000fea4010000000000000000000000000000000000000000003ea401000000000042a40100000000004aa40100000000004ca401000000000054a401000000000056a401000000000058a40100000000005aa4010000000000000000000000000000000000000000004ca401000000000054a401000000000056a401000000000058a4010000000000000000000000000000000000000000002ea601000000000044a601000000000046a60100000000004ea6010000000000000000000000000000000000000000002ea601000000000044a601000000000046a60100000000004ea60100000000000000000000000000000000000000000070a60100000000007aa601000000000082a6010000000000cca60100000000000000000000000000000000000000000070a601000000000074a601000000000082a6010000000000c8a60100000000000000000000000000000000000000000070a601000000000074a601000000000082a6010000000000c8a60100000000000000000000000000000000000000000038a70100000000004ea701000000000054a701000000000058a70100000000000000000000000000000000000000000038a70100000000004ea701000000000054a701000000000058a70100000000000000000000000000000000000000000050a701000000000054a70100000000005aa70100000000005ca70100000000000000000000000000000000000000000072a701000000000076a70100000000007ea701000000000080a701000000000088a70100000000008aa70100000000008ca701000000000090a70100000000000000000000000000000000000000000080a701000000000088a70100000000008aa70100000000008ca701000000000000000000000000000000000000000000a4a7010000000000a8a7010000000000aea7010000000000b0a7010000000000b8a7010000000000baa7010000000000bca7010000000000bea701000000000000000000000000000000000000000000b0a7010000000000b8a7010000000000baa7010000000000bca701000000000000000000000000000000000000000000c0a7010000000000c2a7010000000000cca7010000000000cea7010000000000d6a7010000000000d8a7010000000000daa7010000000000dca701000000000000000000000000000000000000000000cea7010000000000d6a7010000000000d8a7010000000000daa70100000000000000000000000000000000000000000046a801000000000048a80100000000008ca801000000000090a801000000000092a801000000000098a80100000000000000000000000000000000000000000050a801000000000058a80100000000005aa80100000000005ea801000000000060a801000000000066a801000000000068a801000000000078a80100000000007aa80100000000007ca801000000000080a80100000000008ca80100000000000000000000000000000000000000000098a8010000000000b0a8010000000000b2a8010000000000b4a8010000000000c0a8010000000000c2a8010000000000c4a8010000000000c8a801000000000000000000000000000000000000000000e2a8010000000000e8a8010000000000eca8010000000000f2a801000000000018a90100000000004aa9010000000000000000000000000000000000000000006ea901000000000076a901000000000088a90100000000008ca9010000000000000000000000000000000000000000006ea901000000000076a901000000000088a90100000000008ca9010000000000000000000000000000000000000000006ea901000000000072a901000000000088a90100000000008ca901000000000000000000000000000000000000000000caa9010000000000d2a9010000000000d6a9010000000000dea901000000000000000000000000000000000000000000e4a90100000000000eaa0100000000008eaa0100000000009eaa01000000000000000000000000000000000000000000e4a90100000000000eaa0100000000008eaa0100000000009eaa0100000000000000000000000000000000000000000020aa0100000000002eaa01000000000032aa0100000000008caa01000000000000000000000000000000000000000000a2aa010000000000c0aa010000000000deaa010000000000e8aa01000000000000000000000000000000000000000000a2aa010000000000c0aa010000000000deaa010000000000e8aa01000000000000000000000000000000000000000000ecaa010000000000f2aa010000000000f8aa010000000000fcaa01000000000000ab01000000000004ab01000000000000000000000000000000000000000000ecaa010000000000f2aa010000000000f8aa010000000000fcaa01000000000000ab01000000000004ab0100000000000000000000000000000000000000000076ab010000000000ccab010000000000d2ab010000000000e0ab0100000000000000000000000000000000000000000086ab01000000000088ab0100000000009eab010000000000a2ab01000000000000000000000000000000000000000000acab010000000000b6ab010000000000d2ab010000000000e0ab01000000000000000000000000000000000000000000acab010000000000b6ab010000000000d2ab010000000000e0ab01000000000000000000000000000000000000000000acab010000000000b6ab010000000000d2ab010000000000e0ab0100000000000000000000000000000000000000000026ac0100000000003eac0100000000005eac0100000000003aad0100000000000000000000000000000000000000000026ac0100000000003eac0100000000005eac0100000000003aad010000000000000000000000000000000000000000003eac0100000000004cac0100000000006aad0100000000006ead010000000000000000000000000000000000000000003eac0100000000004cac0100000000006aad0100000000006ead010000000000000000000000000000000000000000003eac0100000000004cac0100000000006aad0100000000006ead010000000000000000000000000000000000000000003eac0100000000004cac0100000000006aad0100000000006ead01000000000000000000000000000000000000000000aaad010000000000aead010000000000b6ad010000000000bcad010000000000d8ad010000000000dead01000000000000000000000000000000000000000000a2ae010000000000a6ae010000000000aeae010000000000b4ae010000000000d0ae010000000000d6ae0100000000000000000000000000000000000000000098af0100000000009aaf010000000000a6af01000000000084b001000000000000000000000000000000000000000000aaaf010000000000aeaf010000000000b2af010000000000b6af01000000000000000000000000000000000000000000aaaf010000000000aeaf010000000000b2af010000000000b6af01000000000000000000000000000000000000000000f4af010000000000feaf01000000000000b001000000000004b00100000000000000000000000000000000000000000012b001000000000016b00100000000001cb00100000000005ab00100000000005eb001000000000068b00100000000000000000000000000000000000000000012b001000000000016b00100000000001cb00100000000005ab00100000000005eb001000000000068b001000000000000000000000000000000000000000000b4b0010000000000c6b0010000000000deb0010000000000a2b101000000000000000000000000000000000000000000bcb0010000000000beb0010000000000deb0010000000000a2b101000000000000000000000000000000000000000000e2b0010000000000e6b0010000000000eab0010000000000eeb001000000000000000000000000000000000000000000e2b0010000000000e6b0010000000000eab0010000000000eeb00100000000000000000000000000000000000000000032b101000000000036b10100000000003cb101000000000084b10100000000000000000000000000000000000000000032b101000000000036b10100000000003cb101000000000084b1010000000000000000000000000000000000000000004eb2010000000000a6b2010000000000acb2010000000000bab20100000000000000000000000000000000000000000062b201000000000064b201000000000078b20100000000007cb20100000000000000000000000000000000000000000086b201000000000090b2010000000000acb2010000000000bab20100000000000000000000000000000000000000000086b201000000000090b2010000000000acb2010000000000bab20100000000000000000000000000000000000000000086b201000000000090b2010000000000acb2010000000000bab201000000000000000000000000000000000000000000c0b201000000000018b30100000000001eb30100000000002cb301000000000000000000000000000000000000000000d4b2010000000000d6b2010000000000eab2010000000000eeb201000000000000000000000000000000000000000000f8b201000000000002b30100000000001eb30100000000002cb301000000000000000000000000000000000000000000f8b201000000000002b30100000000001eb30100000000002cb301000000000000000000000000000000000000000000f8b201000000000002b30100000000001eb30100000000002cb3010000000000000000000000000000000000000000004cb30100000000004eb301000000000050b3010000000000d8b3010000000000000000000000000000000000000000004cb30100000000004eb301000000000050b30100000000006cb3010000000000000000000000000000000000000000004cb30100000000004eb301000000000050b301000000000060b301000000000000000000000000000000000000000000eab301000000000040b401000000000046b401000000000054b401000000000000000000000000000000000000000000fab3010000000000fcb301000000000012b401000000000016b40100000000000000000000000000000000000000000020b40100000000002ab401000000000046b401000000000054b40100000000000000000000000000000000000000000020b40100000000002ab401000000000046b401000000000054b40100000000000000000000000000000000000000000020b40100000000002ab401000000000046b401000000000054b4010000000000000000000000000000000000000000009ca2010000000000a0a2010000000000a0a2010000000000aea2010000000000aea2010000000000b0a2010000000000b0a2010000000000f2a3010000000000f2a3010000000000d6a5010000000000d6a50100000000002ca60100000000002ca6010000000000a4a9010000000000a4a9010000000000b2a9010000000000b2a901000000000030ab01000000000030ab01000000000042ab01000000000042ab01000000000054ab01000000000054ab01000000000062ab01000000000062ab01000000000070ab01000000000070ab010000000000e0ab010000000000e0ab0100000000009cad0100000000009cad01000000000050ae01000000000050ae01000000000088ae01000000000088ae01000000000092ae01000000000092ae01000000000048af01000000000048af01000000000082af01000000000082af010000000000a2b0010000000000a2b0010000000000a2b1010000000000a2b10100000000003ab20100000000003ab201000000000048b201000000000048b2010000000000bab2010000000000bab20100000000002cb30100000000002cb301000000000042b301000000000042b3010000000000e4b3010000000000e4b301000000000054b4010000000000000000000000000000000000000000007261775f7665630073747200636f756e74005f5a4e34636f726535736c6963653469746572313349746572244c542454244754243134706f73745f696e635f73746172743137683231633736663939343638653065646545007b636c6f7375726523307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e005f5a4e34636f726533707472347265616431376831626239643039646638396234373532450077726974653c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e007b696d706c2335347d00616476616e63655f62793c636f72653a3a7374723a3a697465723a3a43686172496e64696365733e006e657874005f5a4e34636f726533737472367472616974733131305f244c5424696d706c2475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c5424737472244754242475323024666f722475323024636f72652e2e6f70732e2e72616e67652e2e52616e6765546f244c54247573697a652447542424475424336765743137683633326532303137643665353735396645006e6578743c5b7573697a653b20345d3e00636f6e7461696e735f6e6f6e5f636f6e74696e756174696f6e5f62797465006275696c64657273005f5a4e3131305f244c5424636f72652e2e6f70732e2e72616e67652e2e52616e676546726f6d244c54247573697a6524475424247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c54242475356224542475356424244754242447542435696e6465783137686163396536316662616530626263376145005f5a4e34636f726533666d7439466f726d617474657231327061645f696e74656772616c3137686238656639343965396131613633346545005f5a4e36335f244c5424636f72652e2e63656c6c2e2e426f72726f774d75744572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683636336332373865383138373636393045005f5a4e34636f726533666d74336e756d35335f244c5424696d706c2475323024636f72652e2e666d742e2e55707065724865782475323024666f7224753230246936342447542433666d743137683464336136353331313038303933376445005f5a4e34636f726533666d7439466f726d617474657239616c7465726e617465313768333537326537646636323036356664374500696e646578005f5a4e34636f7265366f7074696f6e31354f7074696f6e244c5424542447542439756e777261705f6f72313768343165333439646137383638346138334500616c69676e5f6f66667365743c75383e005f5a4e34636f72653373747232315f244c5424696d706c24753230247374722447542439656e64735f776974683137683139626662313333653233336465306145005f5a4e34636f726535736c69636532395f244c5424696d706c2475323024247535622454247535642424475424336765743137683233646638653962656438656665346645005f5a4e34636f726533666d74386275696c64657273313044656275675475706c65356669656c6432385f24753762242475376224636c6f7375726524753764242475376424313768636364396362623165623562613563364500656e74727900666d745f696e743c636f72653a3a666d743a3a6e756d3a3a55707065724865782c2075383e005f5a4e34636f726536726573756c743133756e777261705f6661696c65643137683030653934303161326339653536633045005f5a4e34636f726533666d74386275696c6465727338446562756753657435656e7472793137686531623638303262326163636539656445007074720070616464696e670077726974653c636861723e0069735f736f6d653c7573697a653e00676574005f5a4e37355f244c54247573697a65247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c542424753562245424753564242447542424475424336765743137683362336666656535366439303731313345005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243873706c69745f61743137683461343239666364306233623563343945005f5a4e3131305f244c5424636f72652e2e697465722e2e61646170746572732e2e656e756d65726174652e2e456e756d6572617465244c54244924475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e65787431376831623734616564656639323065303665450063686172005f5a4e34636f7265366f7074696f6e31354f7074696f6e244c5424542447542436696e736572743137686265366237313331636461646331646245005f5a4e34636f726536726573756c743139526573756c74244c542454244324452447542438616e645f7468656e3137683138643933303364393238646565393245005f5a4e34636f726536726573756c743139526573756c74244c542454244324452447542438616e645f7468656e313768316532623263316238653933626561654500636f70795f66726f6d5f736c696365007b696d706c2332397d007b696d706c233232357d005f5a4e34636f726533666d7439466f726d6174746572323564656275675f7475706c655f6669656c64315f66696e6973683137683963326264643732306464613133376545007b696d706c2336357d005f5a4e3130385f244c5424636f72652e2e697465722e2e61646170746572732e2e66696c7465722e2e46696c746572244c5424492443245024475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722447542435636f756e743137683631323362313132363938303130326445005f5a4e34636f72653370747235777269746531376830336462313664353065636536366165450072616e6765006f7074696f6e005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f72336e74683137683635613666633036633265613031396645005f5a4e34636f72653373747235636f756e743134646f5f636f756e745f6368617273313768653066306166323562653730356463664500616c69676e5f746f5f6f6666736574733c75382c207573697a653e005f5a4e34636f726533636d70336d696e3137683961303232643031326665326338333745007b696d706c23317d005f5a4e34636f726533666d743372756e313768666639613633333362396633663061614500676574636f756e7400697465725f6d75743c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e006272616e63683c28292c20636f72653a3a666d743a3a4572726f723e007b696d706c2332357d005f5a4e34636f7265336f70733866756e6374696f6e36466e4f6e63653963616c6c5f6f6e63653137683331326365396462383432326365623645005f5a4e34636f726533666d74386275696c64657273313044656275675475706c65356669656c643137686134393061356537663734366534656245005f5a4e34636f72653130696e7472696e736963733139636f70795f6e6f6e6f7665726c617070696e673137683165326664363834393232323263326345005f5a4e34636f726533666d7439466f726d6174746572397369676e5f706c75733137683765363563323535316433616561343445007369676e5f706c7573005f5a4e34636f72653373747235636f756e743233636861725f636f756e745f67656e6572616c5f6361736531376864313333363866323830386530613030450076616c69646174696f6e73005f5a4e34636f726535736c696365346974657238375f244c5424696d706c2475323024636f72652e2e697465722e2e7472616974732e2e636f6c6c6563742e2e496e746f4974657261746f722475323024666f7224753230242452462424753562245424753564242447542439696e746f5f697465723137683765326332623733366531386264656545005f5a4e34636f726533707472376d75745f70747233315f244c5424696d706c2475323024244250246d75742475323024542447542433616464313768333939313037663564323335643062374500497465724d75740047656e657269635261646978006e6578745f696e636c75736976653c636861723e005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243132616c69676e5f6f66667365743137686265366661383332613635626436303545007b696d706c2335337d0064726f705f696e5f706c6163653c26636f72653a3a697465723a3a61646170746572733a3a636f706965643a3a436f706965643c636f72653a3a736c6963653a3a697465723a3a497465723c75383e3e3e005f5a4e34636f7265337074723133726561645f766f6c6174696c653137683034656338646164326362346562306245006d75745f7074720073756d005f5a4e34636f726533666d7439466f726d61747465723770616464696e67313768386664646163386139653836623737364500636d7000696d706c73005f5a4e34636f72653373747232315f244c5424696d706c247532302473747224475424313669735f636861725f626f756e646172793137683034353265303532643135616334353245005f5a4e37355f244c54247573697a65247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c542424753562245424753564242447542424475424336765743137686337356165633633323166633531643545005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542439656e64735f77697468313768383363653331633938643238356662364500696e736572743c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e005f5a4e34636f726533666d74386275696c6465727331304465627567496e6e65723969735f7072657474793137683430666266303734623763353466303545007b696d706c2334317d005f5a4e34636f72653970616e69636b696e673970616e69635f666d743137686436616161656662346334646538633945005f5a4e34636f72653373747235636f756e743131636f756e745f63686172733137683362393037393633646461313835376345007265706c6163653c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e005f5a4e34636f7265366f7074696f6e31354f7074696f6e244c542454244754243769735f736f6d653137686166353061376333383437653666373645006e74683c636f72653a3a7374723a3a697465723a3a43686172496e64696365733e005f5a4e34636f726533737472313176616c69646174696f6e733135757466385f66697273745f627974653137683962396637633933306431356335663945005f5a4e34636f726533666d7438676574636f756e743137683639663830313763343363306364653245005f5a4e34636f72653970616e69636b696e673970616e69635f7374723137683666303932373830653338346562353045005f5a4e34636f726535736c696365366d656d6368723138636f6e7461696e735f7a65726f5f6279746531376861303536386565313833303061353732450072656d00666d745f696e743c636f72653a3a666d743a3a6e756d3a3a4c6f7765724865782c2075383e005f5a4e34355f244c5424244c502424525024247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d74313768613430323766643039663261636331324500666d743c28293e005f5a4e36375f244c5424636f72652e2e61727261792e2e54727946726f6d536c6963654572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d74313768353264643636336235383463633535664500636f70795f6e6f6e6f7665726c617070696e673c75383e00616363756d007b696d706c2334387d007b636c6f7375726523307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542434697465723137686266616536663139613561623764656445006765745f756e636865636b65643c636f72653a3a666d743a3a72743a3a417267756d656e742c207573697a653e006765743c267374723e0070616e69635f646973706c61793c267374723e00756e777261705f6661696c6564002f72757374632f32663662633564323539653761623235646466646433336465353362383932373730323138393138007274005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f7234666f6c64313768623061333862663336373733633236364500636f756e743c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e005f5a4e34636f726533707472347265616431376831653634383335653639376533366630450073756d5f62797465735f696e5f7573697a65005f5a4e34636f726533666d7432727438417267756d656e743861735f7573697a653137686437613231613332353662616362386245005f5a4e3131305f244c5424636f72652e2e697465722e2e61646170746572732e2e656e756d65726174652e2e456e756d6572617465244c54244924475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e657874313768633030313137313163643937383139624500726573756c74005f5a4e37335f244c5424636f72652e2e666d742e2e6e756d2e2e4c6f776572486578247532302461732475323024636f72652e2e666d742e2e6e756d2e2e47656e657269635261646978244754243564696769743137686634306237613733623764393162653445004d61796265556e696e6974007b696d706c2336347d005f5a4e37335f244c54242475356224412475356424247532302461732475323024636f72652e2e736c6963652e2e636d702e2e536c6963655061727469616c4571244c542442244754242447542435657175616c3137686637383434376536346661643333376145005f5a4e3130365f244c5424636f72652e2e6f70732e2e72616e67652e2e52616e6765244c54247573697a6524475424247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c542424753562245424753564242447542424475424336765743137683761383664333261616263343034303345005f5a4e34636f72653463686172376d6574686f647332325f244c5424696d706c247532302463686172244754243131656e636f64655f757466383137683661333732316366346263313738623645005f5a4e34636f726533666d74336e756d313247656e65726963526164697837666d745f696e743137686363663535643038613665313532386645005f5a4e34636f726533666d74336e756d33696d7037666d745f7536343137683238366534643532373433386334363745005f5a4e34636f72653970616e69636b696e673570616e69633137686437373538656430613265383739363145006c6962726172792f636f72652f7372632f6c69622e72732f402f636f72652e353431663036343835316338633866372d6367752e3000726561645f766f6c6174696c653c7573697a653e005f5a4e3130385f244c5424636f72652e2e697465722e2e61646170746572732e2e66696c7465722e2e46696c746572244c5424492443245024475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722447542435636f756e7438746f5f7573697a6532385f24753762242475376224636c6f73757265247537642424753764243137686532646263323632336436376436643345005f5a4e34636f726533666d743131506f737450616464696e673577726974653137683130373832303864313037663934393045006164643c7573697a653e005f5a4e34636f726533666d7439466f726d61747465723977726974655f737472313768353330393765363135313339346565644500696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e2c20636f72653a3a6f70733a3a72616e67653a3a52616e676546726f6d3c7573697a653e3e007b696d706c2331357d00656e64735f776974683c75383e005f5a4e34636f726535736c696365366d656d636872366d656d6368723137683838333063653264646237323666636245006c656e5f75746638005f5a4e34636f72653463686172376d6574686f64733135656e636f64655f757466385f7261773137686230336466376165346464366562316445005f5a4e34636f726533666d74355772697465313077726974655f63686172313768666466623438666364333637346132384500616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23347d3a3a6669656c643a3a7b636c6f737572655f656e7623307d3e00636f7265005f5a4e34636f726533636d7035696d706c7335375f244c5424696d706c2475323024636f72652e2e636d702e2e5061727469616c4f72642475323024666f7224753230247573697a6524475424326c74313768383563303932356636663163316566654500646f5f636f756e745f6368617273005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542431336765745f756e636865636b656431376838333832313033623533356331333034450063656c6c006765743c75382c20636f72653a3a6f70733a3a72616e67653a3a52616e67653c7573697a653e3e004465627567496e6e65720066696e697368005f5a4e34636f726533666d74336e756d313247656e65726963526164697837666d745f696e7431376835383366363662653034373931303631450077726974655f70726566697800636861725f636f756e745f67656e6572616c5f6361736500706f73745f696e635f73746172743c75383e007265706c6163653c636861723e00506f737450616464696e6700697465723c75383e005f5a4e38375f244c5424636f72652e2e7374722e2e697465722e2e43686172496e6469636573247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683862646365633661316137393933386345005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542433676574313768396431656137353833353464396166364500656e756d6572617465005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683563636236663439653430616432356245005f5a4e34636f726535736c69636534697465723136497465724d7574244c54245424475424336e65773137683131393134666634646337396132326545006469676974005f5a4e34636f726535736c69636533636d7038315f244c5424696d706c2475323024636f72652e2e636d702e2e5061727469616c4571244c54242475356224422475356424244754242475323024666f7224753230242475356224412475356424244754243265713137683331383339323064643563373930336445006d656d6368725f616c69676e656400777261705f6275663c636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23317d3a3a777261703a3a7b636c6f737572655f656e7623307d3e005f5a4e34636f726533666d74386275696c6465727331305061644164617074657234777261703137686630613261643433323636313138356545005f5a4e34636f726533666d74386275696c64657273313044656275675475706c653666696e6973683137683262326465366164386361323965353845006974657200666f6c643c7573697a652c20636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c207573697a652c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e005f5a4e34636f72653373747235636f756e743233636861725f636f756e745f67656e6572616c5f6361736532385f24753762242475376224636c6f73757265247537642424753764243137686238333838383631636166343538396545007b636c6f7375726523307d3c2675382c207573697a652c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e00737065635f6e6578743c7573697a653e005f5a4e34636f726534697465723572616e67653130315f244c5424696d706c2475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722475323024666f722475323024636f72652e2e6f70732e2e72616e67652e2e52616e6765244c5424412447542424475424346e6578743137683166316635393732633862353338396245005f5a4e34636f726533737472313176616c69646174696f6e733138757466385f6163635f636f6e745f62797465313768386431353839303565613233346333334500757466385f6163635f636f6e745f62797465006164643c5b7573697a653b20345d3e006e65773c5b7573697a653b20345d3e005f5a4e34636f726535736c6963653469746572313349746572244c542454244754243134706f73745f696e635f73746172743137686632323465323937613136633263656145006e6578743c636f72653a3a736c6963653a3a697465723a3a497465723c636f72653a3a666d743a3a72743a3a417267756d656e743e3e005f5a4e34636f726535617272617938355f244c5424696d706c2475323024636f72652e2e6f70732e2e696e6465782e2e496e646578244c542449244754242475323024666f722475323024247535622454247533622424753230244e24753564242447542435696e6465783137683663646534633833393961376530333445007b696d706c23397d0064656275675f7475706c655f6e6577005f5a4e34636f726533666d74386275696c64657273313044656275675475706c653666696e69736832385f24753762242475376224636c6f737572652475376424247537642431376861393666623161373161643166373535450064656275675f7475706c655f6669656c64315f66696e697368006164643c75383e007b696d706c233138317d00666f6c643c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a6d61703a3a6d61705f666f6c643a3a7b636c6f737572655f656e7623307d3c2675382c207573697a652c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e3e005f5a4e34636f726535736c69636532395f244c5424696d706c2475323024247535622454247535642424475424313873706c69745f61745f756e636865636b65643137683765396534313435376636393734393145006e6578743c636f72653a3a736c6963653a3a697465723a3a497465723c636f72653a3a666d743a3a72743a3a506c616365686f6c6465723e3e007b696d706c2331377d005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542438697465725f6d75743137683030376635633136366631613761373245006172726179005f5a4e34636f7265337374723469746572323253706c6974496e7465726e616c244c5424502447542431346e6578745f696e636c75736976653137683938613230353930343932666138366445005f5a4e35325f244c542463686172247532302461732475323024636f72652e2e7374722e2e7061747465726e2e2e5061747465726e24475424313269735f7375666669785f6f663137683866653837336364343736333664316445005f5a4e34636f726533666d7439466f726d617474657238777261705f6275663137686636336162363038633262616362303045005f5a4e34636f726533666d74336e756d35325f244c5424696d706c2475323024636f72652e2e666d742e2e55707065724865782475323024666f72247532302469382447542433666d743137683438643832613435336137306166353745007b636c6f7375726523307d0070616e69636b696e67005f5a4e35365f244c54247573697a65247532302461732475323024636f72652e2e697465722e2e7472616974732e2e616363756d2e2e53756d244754243373756d3137683739356164323965353439386433333445005f5a4e34636f72653373747232315f244c5424696d706c2475323024737472244754243132636861725f696e64696365733137686466343535663065643137623532303045006765743c75382c207573697a653e005f5a4e34636f7265337074723132616c69676e5f6f66667365743137683534623332333739346162326331313545005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243961735f6368756e6b7331376831643562356538303063366463326238450061735f6368756e6b733c7573697a652c20343e005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e737424753230245424475424336164643137683566666465653639383065666566633145006765745f756e636865636b65643c636f72653a3a666d743a3a72743a3a417267756d656e743e0064656275675f737472756374007b696d706c2332387d0065713c5b75385d2c205b75385d3e0044656275675475706c6500666d745f696e743c636f72653a3a666d743a3a6e756d3a3a55707065724865782c207536343e00636c616e67204c4c564d202872757374632076657273696f6e20312e37312e302d6e696768746c79202832663662633564323520323032332d30352d30392929006974657261746f72005f5a4e34636f726533737472313176616c69646174696f6e7331356e6578745f636f64655f706f696e74313768656364656330303032323838613566354500757466385f66697273745f627974650069735f636861725f626f756e64617279006d696e3c7573697a653e005f5a4e34636f72653373747235636f756e743330636f6e7461696e735f6e6f6e5f636f6e74696e756174696f6e5f627974653137686530636638653465356130663030393045005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137686134633765313364663063343439373145005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243361646431376833356564316564666234363437623138450077726974655f737472005f5a4e34636f726533666d74336e756d313247656e65726963526164697837666d745f696e743137686162643431393537653230363731373445006d617962655f756e696e697400696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e2c20636f72653a3a6f70733a3a72616e67653a3a52616e676546726f6d3c7573697a653e2c203132383e005f5a4e39395f244c5424636f72652e2e7374722e2e697465722e2e53706c6974496e636c7573697665244c54245024475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683536356238663563313134366339666645005f5a4e38315f244c5424636f72652e2e7374722e2e7061747465726e2e2e436861725365617263686572247532302461732475323024636f72652e2e7374722e2e7061747465726e2e2e53656172636865722447542431306e6578745f6d617463683137686231353436643361613035653433333145005f5a4e34636f72653463686172376d6574686f6473386c656e5f75746638313768343935363635353564666635366333654500656e636f64655f757466385f726177006172697468005f5a4e34345f244c54247538247532302461732475323024636f72652e2e6f70732e2e61726974682e2e52656d244754243372656d313768653539336133626230353330333763654500616c6c6f6300747261697473005f5a4e34636f726535736c6963653469746572313349746572244c54245424475424336e65773137683436326338393130346236666239373745005f5a4e34636f7265336e756d32335f244c5424696d706c24753230247573697a652447542431327772617070696e675f6d756c3137683933396664623563663661656266303945006e6577006d656d6368720077726170005f5a4e34636f726533666d74386275696c6465727331304465627567496e6e657235656e7472793137686361303935346134373764373230616545005f5a4e34636f726533666d74386275696c6465727331304465627567496e6e657235656e74727932385f24753762242475376224636c6f73757265247537642424753764243137686336663430636230393339663733626645005f5a4e34636f726533666d74336e756d313247656e65726963526164697837666d745f696e743137683330323730653937613764383866626145007061640070616e6963005f5a4e34636f726533666d74336e756d35335f244c5424696d706c2475323024636f72652e2e666d742e2e4c6f7765724865782475323024666f7224753230246936342447542433666d74313768663235653065383534373535336437314500696d7000616c7465726e617465006d6170005f5a4e3130325f244c5424636f72652e2e697465722e2e61646170746572732e2e6d61702e2e4d6170244c5424492443244624475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722447542434666f6c643137683439653563633739303661396231626645007772697465007b696d706c23377d006d696e5f62793c7573697a652c20666e28267573697a652c20267573697a6529202d3e20636f72653a3a636d703a3a4f72646572696e673e006765743c267374722c207573697a653e005f5a4e34636f726535736c69636535696e64657837345f244c5424696d706c2475323024636f72652e2e6f70732e2e696e6465782e2e496e646578244c542449244754242475323024666f72247532302424753562245424753564242447542435696e64657831376835623336343435386238326632343635450053706c6974496e7465726e616c006e6578743c636861723e0057726974650077726974655f636861723c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e007b696d706c2332367d005f5a4e34325f244c54242452462454247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d74313768633230363132656137383639386165344500666d74007b696d706c23307d004f7074696f6e007b696d706c23387d005f5a4e34636f726533707472376d75745f70747233315f244c5424696d706c2475323024244250246d757424753230245424475424336164643137686433383935323761353331303836366545006765745f756e636865636b65643c267374723e005f5a4e34636f726533666d7439466f726d6174746572313264656275675f73747275637431376838333134343030643138313466376534450070616e69635f737472005f5a4e34636f726533666d74386275696c64657273313564656275675f7475706c655f6e65773137683134383664383033383865636636373745005553495a455f4d41524b455200736c696365005f5a4e34636f7265336d656d377265706c6163653137683665313530623565366261663964346545007061645f696e74656772616c006765743c75383e005f5a4e34636f726535736c6963653469746572313349746572244c54245424475424336e65773137686231373834333338323430613463363745007b696d706c2331397d006e6578745f6d61746368005f5a4e34636f726536726573756c743139526573756c74244c542454244324452447542438616e645f7468656e3137686639613762303833656534636237383245005f5a4e37335f244c5424636f72652e2e666d742e2e6e756d2e2e5570706572486578247532302461732475323024636f72652e2e666d742e2e6e756d2e2e47656e657269635261646978244754243564696769743137683933663339316566393536306361643245005f5a4e34636f72653370747231303264726f705f696e5f706c616365244c542424524624636f72652e2e697465722e2e61646170746572732e2e636f706965642e2e436f70696564244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c542475382447542424475424244754243137683465633534623435323134663763393045005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683334323336653433336537396333623345006c74006368617273005f5a4e34636f72653373747232315f244c5424696d706c247532302473747224475424336765743137686361316261643162613538333362626645006765743c636f72653a3a6f70733a3a72616e67653a3a52616e6765546f3c7573697a653e3e00706f73745f696e635f73746172743c7573697a653e005f5a4e37355f244c54247573697a65247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c54242475356224542475356424244754242447542431336765745f756e636865636b65643137686630663432666234656339376261626145006164643c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e006d6574686f6473005f5a4e34636f726533666d74386275696c64657273313050616441646170746572347772617032385f24753762242475376224636c6f737572652475376424247537642431376862353032353031383864353564626337450063617061636974795f6f766572666c6f7700666d745f753634005f5a4e36385f244c5424636f72652e2e666d742e2e6275696c646572732e2e50616441646170746572247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f7374723137686539366438303337316562386433343445005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243361646431376836343831303738333031643161616237450049746572005f5a4e34636f72653373747232315f244c5424696d706c2475323024737472244754243563686172733137683635643537336338666664393434333645005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f723130616476616e63655f62793137683837343136383366376333383664636245006e6578745f636f64655f706f696e743c636f72653a3a736c6963653a3a697465723a3a497465723c75383e3e005f5a4e39335f244c5424636f72652e2e736c6963652e2e697465722e2e4368756e6b73244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137686264343939663734373230663065386245004f7264006164643c267374723e007b696d706c23367d00616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23357d3a3a656e7472793a3a7b636c6f737572655f656e7623307d3e004465627567536574005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f666d743137683565373464633863623261616161323645007b696d706c23327d005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542434697465723137686331616261316236653465646465623545005f5a4e34636f726533666d7439466f726d6174746572336e65773137686165623034366666366431666231663445005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243361646431376838353436653232346135313966363633450064656275675f7374727563745f6e657700746f5f7538005f5a4e34636f726533636d7035696d706c7336395f244c5424696d706c2475323024636f72652e2e636d702e2e5061727469616c4571244c54242452462442244754242475323024666f7224753230242452462441244754243265713137683436393566636435376362636161326145005f5a4e34636f726533666d743577726974653137683537653362636463656237646630393145006578706563745f6661696c6564006c656e5f6d69736d617463685f6661696c006f707300696e7472696e736963730073756d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e005f5a4e34636f7265336d656d377265706c61636531376838363534306363336630326138396663450069735f6e6f6e653c7573697a653e00697465723c5b7573697a653b20345d3e00696e746f5f697465723c5b7573697a653b20345d3e005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683366313636623661373436326234373945005f5a4e34636f726533666d7432727438417267756d656e7433666d74313768363232636537653835383430326338654500666d745f696e743c636f72653a3a666d743a3a6e756d3a3a4c6f7765724865782c207536343e00657175616c3c75382c2075383e005f5a4e34636f726535736c696365366d656d63687231326d656d6368725f6e616976653137686363623962373463393862393633336245006d656d6368725f6e6169766500616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23347d3a3a66696e6973683a3a7b636c6f737572655f656e7623307d3e00636f6e73745f707472005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f723373756d313768616537613566613764646461346162384500757466385f69735f636f6e745f62797465006e6578743c636f72653a3a666d743a3a72743a3a417267756d656e743e005f5a4e34636f726533666d74386275696c64657273313664656275675f7374727563745f6e65773137686135363836656238343531653037323245005f5a4e34636f72653970616e69636b696e67313370616e69635f646973706c6179313768663965353336303933393038663832624500656e64735f776974683c636861723e0065713c75382c2075383e007b696d706c23347d005f5a4e34636f726533737472313176616c69646174696f6e733137757466385f69735f636f6e745f6279746531376861396331376363326537313134623836450073706c69745f61745f756e636865636b65643c75383e0073706c69745f61743c75383e005f5a4e34636f72653373747235636f756e74313873756d5f62797465735f696e5f7573697a653137683733663965326535343130353136333245006e6578743c636f72653a3a666d743a3a72743a3a506c616365686f6c6465723e00417267756d656e74005f5a4e37355f244c54247573697a65247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c54242475356224542475356424244754242447542431336765745f756e636865636b6564313768656630633435353430343632353962624500636f6e7461696e735f7a65726f5f62797465005f5a4e37395f244c5424636f72652e2e726573756c742e2e526573756c74244c5424542443244524475424247532302461732475323024636f72652e2e6f70732e2e7472795f74726169742e2e54727924475424366272616e63683137683034646133323232663535363066313845005f5a4e34636f7265366f7074696f6e31336578706563745f6661696c65643137686332333330616533386638616564396545005f5a4e34636f726533707472376d75745f70747233315f244c5424696d706c2475323024244250246d7574247532302454244754243361646431376837336363316163653933303039363536450073756d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e2c207573697a653e005f5a4e35365f244c54247573697a65247532302461732475323024636f72652e2e697465722e2e7472616974732e2e616363756d2e2e53756d244754243373756d32385f24753762242475376224636c6f73757265247537642424753764243137683665653564323561643365666465373945007369676e5f61776172655f7a65726f5f70616400726561643c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e006e6578743c7573697a653e00756e777261705f6f723c267374723e005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243136616c69676e5f746f5f6f6666736574733137683265333033653231353164623038353745005f5a4e34636f726535736c69636532395f244c5424696d706c2475323024247535622454247535642424475424336765743137683037666466393631613031323632356145006e65773c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e007b696d706c2334347d0077726974655f7374723c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e577269746524475424313077726974655f636861723137683239666437616639333939643762333645005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243135636f70795f66726f6d5f736c69636531376c656e5f6d69736d617463685f6661696c3137686531663934356265353831313135613845006c6962726172792f616c6c6f632f7372632f6c69622e72732f402f616c6c6f632e643733613839653266303538366464312d6367752e30004974657261746f7200636f756e745f6368617273005f5a4e34636f72653469746572386164617074657273336d6170386d61705f666f6c6432385f24753762242475376224636c6f73757265247537642424753764243137686265643362346664336632356561633645005f5a4e34636f7265366f7074696f6e31354f7074696f6e244c542454244754243769735f6e6f6e653137683036303537623832613939663564313445005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542438616c69676e5f746f3137686361663565313535373365303734303345007b696d706c2331317d005f5a4e34636f726533636d70366d696e5f62793137683961363365346463336265666132393045005f5a4e34636f7265336d656d31326d617962655f756e696e697432304d61796265556e696e6974244c54245424475424357772697465313768643262633963366561386361383161624500656e636f64655f75746638005f5a4e34636f726533666d743557726974653977726974655f666d743137683364623431343565346436363932376245006669656c64007b696d706c2334307d005f5a4e36305f244c5424636f72652e2e63656c6c2e2e426f72726f774572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137686163386261333334363731373261333845005f5a4e34636f726533666d74336e756d35325f244c5424696d706c2475323024636f72652e2e666d742e2e4c6f7765724865782475323024666f72247532302469382447542433666d743137683039663834613031663936303437366145006e6578743c75383e00746f5f7573697a65006d656d005f5a4e34636f7265337074723577726974653137683934303032343231393363646338316545005f5a4e38395f244c5424636f72652e2e6f70732e2e72616e67652e2e52616e6765244c54245424475424247532302461732475323024636f72652e2e697465722e2e72616e67652e2e52616e67654974657261746f72496d706c2447542439737065635f6e65787431376834303038636235396134653064623339450061735f7573697a65006164643c636f72653a3a666d743a3a72743a3a417267756d656e743e00696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e005f5a4e34636f7265336e756d32335f244c5424696d706c24753230247573697a652447542431327772617070696e675f73756231376838643635306338643866353735643162450069735f70726574747900616461707465727300726561643c636861723e007b696d706c23337d00636861725f696e646963657300616c69676e5f746f3c75382c207573697a653e007772617070696e675f6d756c0077726974653c75383e005f5a4e35305f244c5424753634247532302461732475323024636f72652e2e666d742e2e6e756d2e2e446973706c6179496e742447542435746f5f75383137683636316463333963356464386666653545007061747465726e0069735f7375666669785f6f66005f5a4e34636f726535736c696365366d656d63687231346d656d6368725f616c69676e6564313768643864383232303663636532343531614500526573756c7400506164416461707465720070616e69635f666d74005f5a4e34636f726533666d7439466f726d6174746572337061643137683433336537613934646232626438653245005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f7374723137683865303931326361326264646233386345005f5a4e34636f726533666d7432727431325553495a455f4d41524b455232385f24753762242475376224636c6f7375726524753764242475376424313768643137376134333532613130653633314500466e4f6e6365006e756d005f5a4e38315f244c5424636f72652e2e7374722e2e697465722e2e4368617273247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722447542435636f756e743137686638633866336432633063356164333545005f5a4e34636f726533666d7439466f726d617474657231397369676e5f61776172655f7a65726f5f7061643137683136323439616566366630343733333545006e65773c75383e007b696d706c23357d005f5a4e34636f726533636d70334f7264336d696e31376861623865636338303366663033636364450072756e005f5a4e34636f726533666d74386275696c64657273313044656275675475706c653969735f7072657474793137683131646663373739346165376162303045005f5a4e34636f726533666d7439466f726d617474657231327061645f696e74656772616c313277726974655f70726566697831376838346635386564303837613362643933450066756e6374696f6e00466f726d61747465720066696c746572006d61705f666f6c64005f5a4e38315f244c5424636f72652e2e7374722e2e697465722e2e4368617273247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683064323235303663643135633337363345007b696d706c2337307d005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683634663237353939353136663335636545005f5a4e35355f244c542424524624737472247532302461732475323024636f72652e2e7374722e2e7061747465726e2e2e5061747465726e24475424313269735f7375666669785f6f663137686536396533336230613062663235373545007772617070696e675f7375620077726974655f666d743c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e005f5a4e35616c6c6f63377261775f766563313763617061636974795f6f766572666c6f7731376837363964333737343539393364316265450063616c6c5f6f6e63653c636f72653a3a666d743a3a72743a3a5553495a455f4d41524b45523a3a7b636c6f737572655f656e7623307d2c2028267573697a652c20266d757420636f72653a3a666d743a3a466f726d6174746572293e003a000000020000000000510000003400000063617061636974795f6f766572666c6f77002f0000007261775f766563002a000000616c6c6f630000000000ea1b0000020051000000272600006a01000077726974653c636861723e00322200006d617962655f756e696e697400be2400006272616e63683c28292c20636f72653a3a666d743a3a4572726f723e00e90000006d75745f7074720010230000696e736572743c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e00070400007b696d706c2334317d003d1c0000636f70795f6e6f6e6f7665726c617070696e673c75383e005d060000466f726d617474657200aa2300007b696d706c2331377d001c200000737065635f6e6578743c7573697a653e00c01c0000706f73745f696e635f73746172743c7573697a653e00a71b0000617269746800d8180000446562756753657400091b00007b696d706c2332357d008c240000526573756c7400372100006e6578745f636f64655f706f696e743c636f72653a3a736c6963653a3a697465723a3a497465723c75383e3e0034000000726561645f766f6c6174696c653c7573697a653e00651d0000697465723c5b7573697a653b20345d3e00252200007265706c6163653c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e00dd1f00007b636c6f7375726523307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e00311d000073706c69745f61745f756e636865636b65643c75383e00182200007265706c6163653c636861723e00f622000069735f6e6f6e653c7573697a653e007f1d00006765743c267374722c207573697a653e000c2500007b696d706c2332367d009321000069735f636861725f626f756e64617279006d240000726573756c7400581b000066756e6374696f6e00d31f0000636f756e7400960600007061645f696e74656772616c004b1d0000616c69676e5f746f5f6f6666736574733c75382c207573697a653e00c51d00006c656e5f6d69736d617463685f6661696c00da0000006164643c75383e00a81c00006e65773c75383e00fa030000646967697400211b0000666d743c28293e00c11b000070616e69636b696e670003230000756e777261705f6f723c267374723e00b1200000636f6e7461696e735f6e6f6e5f636f6e74696e756174696f6e5f6279746500cd000000616c69676e5f6f66667365743c75383e00f71c00006e65773c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e000b2400007b696d706c2331397d00962300007772617070696e675f737562006f060000616c7465726e61746500822200006c7400aa1f00006d61705f666f6c6400bd20000073756d5f62797465735f696e5f7573697a6500ae010000417267756d656e7400372200004d61796265556e696e6974009a050000666d7400b11b000072656d001e2300006578706563745f6661696c656400f1020000666d745f696e743c636f72653a3a666d743a3a6e756d3a3a4c6f7765724865782c2075383e000b1f0000636f6e7461696e735f7a65726f5f62797465004f13000072756e00122100007b696d706c2334347d00d82100007b696d706c2332387d003313000077726974655f707265666978005d1b0000466e4f6e6365002a1e00006765743c267374723e005b000000636f6e73745f70747200032200006e6578745f6d6174636800b31d00006765743c75382c20636f72653a3a6f70733a3a72616e67653a3a52616e67653c7573697a653e3e00e5020000666d745f696e743c636f72653a3a666d743a3a6e756d3a3a55707065724865782c2075383e006322000077726974653c75383e00340100006164643c7573697a653e00971c00004974657200dd14000064656275675f7374727563745f6e6577001c1b00007b696d706c2335337d00b30000006164643c636f72653a3a666d743a3a72743a3a417267756d656e743e005920000073747200f81b000070616e69635f646973706c61793c267374723e000a1d0000697465723c75383e00c01d0000636f70795f66726f6d5f736c69636500931f00006d617000d32100007061747465726e00d9020000666d745f696e743c636f72653a3a666d743a3a6e756d3a3a4c6f7765724865782c207536343e005617000066696e69736800f50300007b696d706c2332397d00ab240000616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23347d3a3a66696e6973683a3a7b636c6f737572655f656e7623307d3e0072240000756e777261705f6661696c6564005a1c00006e6578743c75383e00ff20000053706c6974496e7465726e616c008d200000646f5f636f756e745f6368617273008a1c00006e6578743c636f72653a3a666d743a3a72743a3a417267756d656e743e004b1c0000736c696365006a17000044656275675475706c6500d81f0000746f5f7573697a65009c1c0000706f73745f696e635f73746172743c75383e00ca2000006974657200791f000073756d007d2200007b696d706c2335347d00cd1c00007b696d706c2337307d001e1e00006765745f756e636865636b65643c636f72653a3a666d743a3a72743a3a417267756d656e743e009e240000616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23357d3a3a656e7472793a3a7b636c6f737572655f656e7623307d3e00551a00007b696d706c23307d007b200000636861725f636f756e745f67656e6572616c5f6361736500f021000069735f7375666669785f6f66009d1f0000666f6c643c7573697a652c20636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c207573697a652c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e0025120000777261705f6275663c636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23317d3a3a777261703a3a7b636c6f737572655f656e7623307d3e00da1a000077726974655f666d743c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e00e3010000666d745f753634002a000000636f726500581d000061735f6368756e6b733c7573697a652c20343e000813000064656275675f7475706c655f6669656c64315f66696e697368009c0100005553495a455f4d41524b4552008e1f00006164617074657273007c2300007772617070696e675f6d756c007e1f00007b636c6f7375726523307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e009f2100006765743c636f72653a3a6f70733a3a72616e67653a3a52616e6765546f3c7573697a653e3e00a60000006164643c5b7573697a653b20345d3e00c71f0000636f756e743c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e00e51c0000696e746f5f697465723c5b7573697a653b20345d3e002d1f0000666f6c643c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a6d61703a3a6d61705f666f6c643a3a7b636c6f737572655f656e7623307d3c2675382c207573697a652c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e3e00871800007b696d706c23317d00ec2500006368617200bd1f000066696c74657200ed1f0000656e756d657261746500e71e00006d656d6368725f6e6169766500c61b000070616e69635f666d74008906000070616464696e67002e0300007b696d706c2336347d00681f00007b696d706c2334387d008c1800007772617000ca19000064656275675f7475706c655f6e657700e91400007b696d706c23327d00b301000061735f7573697a65006d1f000073756d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e0078220000696d706c7300ac1b00007b696d706c233232357d00631f0000616363756d00d8190000577269746500df1b000070616e6963007e1c00006e6578743c636f72653a3a666d743a3a72743a3a506c616365686f6c6465723e0079210000636861727300531b00006f707300f12500006d6574686f647300c81e000065713c75382c2075383e00172100006e6578743c636861723e00950500007b696d706c2336357d00ac210000656e64735f776974683c636861723e00132200006d656d00eb2100007b696d706c23337d00041c000070616e69635f737472007c1700006669656c6400be2200004f72640097010000727400de010000696d7000f71f00006e6578743c636f72653a3a736c6963653a3a697465723a3a497465723c636f72653a3a666d743a3a72743a3a506c616365686f6c6465723e3e00721c00006e6578743c7573697a653e00f21c0000497465724d75740069130000777269746500991d0000656e64735f776974683c75383e00b118000069735f70726574747900661c00006e6578743c5b7573697a653b20345d3e009f1800004465627567496e6e657200dd180000656e74727900471f0000616476616e63655f62793c636f72653a3a7374723a3a697465723a3a43686172496e64696365733e00d402000047656e65726963526164697800ba21000074726169747300fd020000666d745f696e743c636f72653a3a666d743a3a6e756d3a3a55707065724865782c207536343e005a1a000077726974655f7374723c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e00f22000006e657874003a1f000073756d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e2c207573697a653e003e1700007b696d706c23347d00ee14000077726974655f73747200f62500006c656e5f7574663800a222000065713c5b75385d2c205b75385d3e005d010000726561643c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e003e1d000073706c69745f61743c75383e00042100006e6578745f696e636c75736976653c636861723e001c0300007b696d706c2331317d0050010000726561643c636861723e007f09000070616400af1f00007b636c6f7375726523307d3c2675382c207573697a652c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e00731a000077726974655f636861723c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e0043210000757466385f66697273745f6279746500bf1800007b696d706c23357d00032000006e6578743c636f72653a3a736c6963653a3a697465723a3a497465723c636f72653a3a666d743a3a72743a3a417267756d656e743e3e00b12200006d696e5f62793c7573697a652c20666e28267573697a652c20267573697a6529202d3e20636f72653a3a636d703a3a4f72646572696e673e00ff1100006e657700652300006e756d007701000077726974653c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e00081e0000696e64657800e42200004f7074696f6e00e922000069735f736f6d653c7573697a653e00d81400006275696c646572730086210000636861725f696e646963657300a523000063656c6c00c00000006164643c267374723e00171d00006765743c75382c207573697a653e00431e00007b696d706c23367d00911e00006765743c75383e005b1700007b636c6f7375726523307d002b210000757466385f69735f636f6e745f6279746500281f00004974657261746f7200621b000063616c6c5f6f6e63653c636f72653a3a666d743a3a72743a3a5553495a455f4d41524b45523a3a7b636c6f737572655f656e7623307d2c2028267573697a652c20266d757420636f72653a3a666d743a3a466f726d6174746572293e00f31e00006d656d6368725f616c69676e656400241d0000616c69676e5f746f3c75382c207573697a653e00721d00006765745f756e636865636b65643c636f72653a3a666d743a3a72743a3a417267756d656e742c207573697a653e00410100006164643c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e00fa1d0000697465725f6d75743c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e00df2200006f7074696f6e0003260000656e636f64655f757466385f726177002621000076616c69646174696f6e7300a01e0000636d7000c421000067657400361e00006765745f756e636865636b65643c267374723e00291300007b696d706c23377d00551c00007b696d706c233138317d00231f00006974657261746f72001812000064656275675f737472756374007f1e0000696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e2c20636f72653a3a6f70733a3a72616e67653a3a52616e676546726f6d3c7573697a653e3e00541f00006e74683c636f72653a3a7374723a3a697465723a3a43686172496e64696365733e0015260000656e636f64655f7574663800751800005061644164617074657200db1e00006d656d63687200bf2100007b696d706c23387d00111c0000696e7472696e7369637300fe240000696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e2c20636f72653a3a6f70733a3a72616e67653a3a52616e676546726f6d3c7573697a653e2c203132383e001220000072616e676500d22400007b696d706c2331357d007c0600007369676e5f61776172655f7a65726f5f70616400620600007369676e5f706c7573002f000000707472004100000064726f705f696e5f706c6163653c26636f72653a3a697465723a3a61646170746572733a3a636f706965643a3a436f706965643c636f72653a3a736c6963653a3a697465723a3a497465723c75383e3e3e006f200000636f756e745f636861727300b41c00006e65773c5b7573697a653b20345d3e0016130000506f737450616464696e670067210000757466385f6163635f636f6e745f6279746500481e0000696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e00902200007b696d706c23397d005c130000676574636f756e740091240000616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23347d3a3a6669656c643a3a7b636c6f737572655f656e7623307d3e00d12200006d696e3c7573697a653e0021030000746f5f753800ce0400007b696d706c2334307d00aa1e0000657175616c3c75382c2075383e00cd240000617272617900000000000e00000002000000000051000000000000000e0000000200510000002726000000000000412a000000726973637600012000000004100572763634693270305f6d3270305f613270305f633270300058000000040034000000010101fb0e0d0001010101000000010000016c6962726172792f616c6c6f632f73726300007261775f7665632e727300010000000009022465010000000000038a040105050a030109020001090c00000101771e000004005e030000010101fb0e0d0001010101000000010000016c6962726172792f636f72652f7372632f6f7073006c6962726172792f636f72652f7372632f707472006c6962726172792f636f72652f7372632f666d74006c6962726172792f636f72652f737263006c6962726172792f636f72652f7372632f736c6963652f69746572006c6962726172792f636f72652f7372632f697465722f747261697473006c6962726172792f636f72652f7372632f737472006c6962726172792f636f72652f7372632f69746572006c6962726172792f636f72652f7372632f697465722f6164617074657273006c6962726172792f636f72652f7372632f6d656d006c6962726172792f636f72652f7372632f6d6163726f73006c6962726172792f636f72652f7372632f736c696365006c6962726172792f636f72652f7372632f6e756d006c6962726172792f636f72652f7372632f6172726179006c6962726172792f636f72652f7372632f63686172000066756e6374696f6e2e7273000100006d6f642e72730002000072742e72730003000070616e69636b696e672e7273000400006e756d2e727300030000636f6e73745f7074722e727300020000696e7472696e736963732e7273000400006d75745f7074722e7273000200006d6f642e7273000300006d6163726f732e7273000500006974657261746f722e72730006000076616c69646174696f6e732e727300070000616363756d2e727300060000636d702e72730004000072616e67652e7273000800006d61702e72730009000066696c7465722e727300090000636f756e742e727300070000697465722e7273000700006d6f642e7273000a00006f7074696f6e2e7273000400006d6f642e7273000b00006d6f642e727300070000696e6465782e7273000c00007472616974732e7273000700006d6f642e7273000c000075696e745f6d6163726f732e7273000d0000697465722e7273000c0000656e756d65726174652e72730009000063656c6c2e7273000400006275696c646572732e727300030000726573756c742e7273000400006d617962655f756e696e69742e7273000a00006d6f642e7273000e0000636d702e7273000c00007061747465726e2e7273000700006d656d6368722e7273000c00006d6574686f64732e7273000f000061726974682e727300010000000009029ca201000000000003f90101040205090a03860a090000010403050503d375090200010902000001010404000902a0a2010000000000033301050e0a030f09020001090c000001010402000902aea201000000000003ea030105010a0300090000010902000001010405000902b0a201000000000003d2010105170a03130906000106039a7e0918000103e60109040001039a7e0924000105150603e80109020001051e0302090e00010406050d03b505091a00010407050903d20d090200010405051e03fa6c0904000104070509038613090400010406050d03ae72090800010407050903d20d090200010405051503fb6c09080001040705090385130902000106030009040001040505170603f56c0908000106039a7e0906000105140603f901090400010515030209040001051e037f091c000105150302090400010406050d03a305090200010407050903d20d090200010408050d039c73090c00010407050903e40c0902000106038f6b090a000104050514060381020902000105150301090400010408050d038b06090800010405051503f67909020001051e0302090a000105150301090200010406050d039905090400010407050903d20d090200010408050d039c73090c00010407050903e40c0902000106038f6b090800010408050d06038d08090400010405053e03827a09060001050d030209020001050a030109140001060b0300090200010904000001010409000902f2a301000000000003dd090105090a03e003091e0001051303a77c090c000106039b76090c000105090603f70d09040001051303ee7b0904000105190305090200010603967609020001050f0603fb090902000105090603000902000103857609040001040a051806038601090200010603fa7e09040001040b05150603b113090400010408050d03dc7409040001040c0505038c7809020001040a051803ed0009080001040d051c03af7f09020001040a051803d100090200010409050d03e50809020001050f031009020001050906030009020001052306030909020001051a06030009040001050906038d0409040001051a03f97b09020001051b03e90009020001053103a47f09060001051503dc000904000106038d7509060001050606039d0a09200001060b0300091c0001050003e3750904000104020509060394090926000106030009060001040905110603f900090400010402050903cd00090a000106030009040001040905110603b37f090400010603f3750914000105090603800b09020001040e05340353090600010409050d032e090400010603ff740910000105150603f30a090200010530030a0904000105230603000904000105300300090200010383750906000105090603800b090c0001040e0534035309040001040f050c039a7a090200010409050d039406090200010603ff74090c000105240603970a090a00010511030109040001030109140001050903fb7e090e0001040e053403bf01090800010409050d03c27e09080001051103fa00091000010603f175091000010603910a090200010301090400010603ee7509080001040e05340603d30a090200010906000001010409000902d6a501000000000003f2090105140a0301091c0001051103010904000105140302090e0001052c060300090200010b03000912000103897609040001050a0603f80909020001060b0300090a000109040000010104090009022ca601000000000003bb0a01041505120a039b7a090200010409050c03e7050916000104160509039a78090200010409050c03e607090800010518030509040001051d060300090400010406050d0603dc7c09040001040b050903b87b09040001040c05000603a97d09120001041305260603910109040001051106030009020001040b05100603c70109040001040e053403fb0709040001040f050c039a7a09020001040a051803997c09020001040c050d03a07f0904000105080301090800010516030a090400010505035b0904000105110306090400010508032109040001051a0305090400010505035a090400010511060300090200010505030009040001050c06032909040001051e030509040001051203010904000105050351090400010511060300090200010505030009040001050d06032f090400010413050903cb00090200010603f47e09040001040a051806038601091e0001040c050d03a07f090400010508030109040001060359090400010603330908000106034d09040001050c06033b09040001050006034509040001051a060338090400010511035a0904000106030009040001051e06032e09040001051203010904000105050351090400010511060300090600010505030009040001050d06032f090200010413050903cb00090600010417050c03cc000904000105090304090200010418050c037d0904000104170513030f0904000104190509032c090800010603ec7d0904000104150603bc0709020001041903d87a090400010603ec7d0904000104150603bc07090200010603c4780902000104090603d40a0904000105120304090400010412050803c3750908000106036509040001040a051806038601090200010603fa7e09040001040b05150603b113090400010408050d03dc7409040001040c0505038c7809020001040a051803ed0009080001040d051c03af7f09020001040a051803d100090200010402051f03bb0c09040001041a0545036509060001051603800e09080001040a051803e065090600010603fa7e09040001040b05150603b113090200010408050d03dc7409040001040c0505038c7809020001040a051803ed0009080001040d051c03af7f09020001040a051803d100090200010603fa7e090200010386010902000103fa7e09020001040b05150603b113090600010408050d03dc7409040001040c0505038c7809020001040a051803ed0009080001040d051c03af7f09020001040a051803d100090200010603fa7e09020001041205150603c7000922000105000603b97f09060001051b0603fe00090e00010534060300090400010533030009020001051b030009040001041b050d0603e7080902000104120505039a77090400010509035b09020001050c030609020001041c03e80a090200010603b87409020001041a053806039908091200010406050d03867f09040001040a051803e779090600010603fa7e09020001041205190603d0000904000105120301090200010507032309020001050606030009040001051203000902000106035d09020001050503230902000105110360090400010507032009020001050606030009040001051206035d090200010323090200010505060300090200010507030009040001050603000904000105120300090200010505030009020001051206035d0902000105050323090200010511036009020001050703200904000105060603000904000105120300090200010505030009020001040a05180603120904000104120511034e09040001040a05180332090200010603000906000103fa7e090400010386010904000103fa7e09040001038601090600010412051206035d090600010408050d03aa07090200010412050703e7780902000105060603000904000105120300090200010505030009020001040a05180603120904000104120511035e09020001040a05180322090200010603fa7e090400010412051b0603fe00090200010534060300090400010533030009020001051b030009040001041b050d0603e7080902000104120505039a7709040001050d0367090200010409051403f60909020001051b0317090400010535037009060001051503100904000106038d750906000103f30a09260001053006030a0904000105230603000904000105300300090200010383750906000105090603800b090e0001040e0534035309040001040f050c039a7a090200010409050d039406090200010603ff74090c000105280603e30a090a00010515030109040001050903b07e090e0001040e053403bf0109080001040f050c039a7a090400010409050d03a804090400010603eb7609100001040e05340603d30a0902000104090506031609040001060b0300091400010904000001010404000902a4a901000000000003ed000105050a030709020001090c000001010409000902b2a901000000000003b7080105090a03bb7909180001050b03c90609080001050903b77909040001050503c90609080001050e030e09020001040a051803bc78090400010603fa7e0904000103860109040001040905150603cb0709220001051406030009020001051506030109020001052d0603000904000105150300090400010510060313090600010505060300090200010511060301090200010505060300090400010511060301090400010533036f09020001050503110904000105150304090200010505030f090600010403050c039978090600010603ed7e090a0001051d0603960109040001051b0603000902000103ea7e09020001040905090603eb080902000105190301090400010505030e090800010403050c039978090600010603ed7e090a0001051d0603960109040001051b0603000902000103ea7e09020001040905090603ec0809020001052d0307090400010406050d03ac7e090200010403050903eb7909040001051a060300090200010509030009020001040905110603cc0709040001040a051803b078090200010409051d03b90709100001040a051803c778090400010603fa7e0904000103860109080001040905150603bd0709120001051406030009020001051506030109020001052d060300090400010515030009040001040305090603c67809060001051a060300090200010509030009040001040905110603bc0709040001040a051803c078090200010409051a03d707090a00010418050c03fc78090400010603a77e090600010409051a0603dd08090200010418050c03fc78090400010409051a038407090400010406050d03c27e090400010409050903bf0109040001052106030009040001050903000908000103a2770906000105020603e20809060001060b030009100001090400000101041e00090230ab01000000000003ba0501040905090a03ba0609000001091200000101041e00090242ab01000000000003d50501040905090a039f0609000001091200000101042000090254ab01000000000003f10c0105050a030109020001090c00000101041500090262ab010000000000038a0f01040405050a038b7209020001090c00000101040500090270ab010000000000039901010408050d0a03f30609060001040505000603f3770908000106039301090800010421050903d602090200010405051403ea7c090400010603ad7f09080001052306032a0902000103e900090800010603ed7e090400010418050c0603ed03090a00010405050903817d090a0001050e032e09160001060b0300090200010418050d0603d20209040001090e00000101041f000902e0ab010000000000031e010413050c0a03ce0409460001041a0523039c0d091800010423050d03d26e09040001041f034a090a00010301090400010413050c03c704090e00010424051903b17e090800010418050c0342090a00010425050803cb7d09080001050b030d0906000106034809040001050c0603390902000105090304090c0001050b037b090200010402051f03890d09060001051b03010908000104250508039273090400010603ac7f090e000105100603eb00090600010406050d03b406090400010425051503c679090400010529030409060001041b050d03e508090200010425050503c67609020001051503d2000908000105290304090a0001041b050d03e408090200010425050503c67609020001050903db0009080001050b037209020001050c03580906000105090304090c0001050b037b09020001060348090400010603e1000904000106039f7f09040001050c06033909060001050b037f090c000106034809080001042405200603b403090200010511060300090200010418050c0603ac7f090800010423050d03fb7d090200010424051c03dd02090400010603c87c09040001041f051006032109140001051103010906000106035e090e0001041a050906038912090800010603f76d09040001041f050606032a09100001060b0300091a000109040000010104090009029cad01000000000003a20101052b0a0301090c00010426050803f60b09020001050d031f09040001050f0363090800010513032009060001050d06030009040001051206030109080001050d06030009040001050f060361090c00010513032209060001050d06030009040001051206030109080001050d06030009060001051206030109080001050d060300090400010512060303090c0001050d06030009060001051206030109080001050d06030009060001051206030109080001050d06030009060001051206030109080001050d06030009040001040905090603dc73090a000105060301090a0001060b030009020001090400000101040900090250ae01000000000003be010105090a0301090200010506030109300001060b030009020001090400000101040900090288ae01000000000003c5010105090a030109000001090a00000101040900090292ae01000000000003c9010105090a030109020001052b0359090c00010426050803f60b09020001050d031f09040001050f0363090800010513032009060001050d06030009040001051206030109080001050d06030009040001050f060361090c00010513032209060001050d06030009040001051206030109080001050d06030009060001051206030109080001050d060300090400010512060303090c0001050d06030009060001051206030109080001050d06030009060001051206030109080001050d06030009060001051206030109080001050d06030009040001040905090603dc73090a000105060328090a0001060b030009020001090400000101040900090248af01000000000003cd010105090a0301090200010371091e00010506031009140001060b030009020001090400000101041f00090282af01000000000003b3020105170a0301091200010420050903f10709040001041f03a078090200010603ba7d0908000105100603b602090400010409050903c10b09040001041f050006038972090400010409050903f70d09040001041f05100603bf740904000105000603ca7d09020001051e0603c002090400010603c07d0904000105140603b702090a00010409050903be0909040001041f051503c376091600010603c87d09020001040905090603f50b090e0001041f051e03cb76090a00010409050903b50909020001042003a70309040001041f051103a673090200010409051403e406090c00010603da7609040001041f05210603bb02090200010409051703e806090400010415050903f002090800010409051303947d090a0001051403010904000103010904000105180301090800010509037709080001041f0511039c79091400010409050903e40609040001041f0511039c79090a00010409050903b80909080001041f050006038b740912000105090603b502090200010311090400010506030209060001060b030009100001090400000101041f000902a2b001000000000003d3030105170a03a87f091200010420050903aa0709080001041f03d67809020001031209040001050603c90009040001060b03000910000103a97c0904000105100603fd02090400010409050903fa0a09040001041f050006038972090400010409050903f70d09040001041f051006038675090400010514030a090200010409050903ee0809020001041f051503937709180001051103020902000105140374090a00010409050903f70809020001041f0515038a77091800010409051403a706090200010603da7609040001041f052106038203090200010409051703a106090400010415050903f002090800010409051303947d090a0001051403010904000103010904000105180301090800010509037709080001041f051103e379091e00010409050903f108090800010916000001010409000902a2b101000000000003e40f0105090a03907c090c0001041f050503a376090c00010409050903cf0d090c0001041f050c03fd72090e0001050006039c7d09020001050c03e40209040001039c7d09020001042005090603a60a09020001041f051403c07809020001050006039a7d090a0001051403e60209020001040905090603910b09080001041f051403ef740906000104090509038f0909020001041f051503f2760914000104090509038e0909020001041f03f776091600010409050603fd0c09040001060b0300090a0001090400000101041a0009023ab2010000000000038a1a01050d0a030109020001090c00000101040500090248b2010000000000039901010408050d0a03f30609060001040505000603f3770908000106039401090c00010421050903d502090200010405051403ea7c090400010427052d03ef03090800010405052303d27c090800010603ec7e090400010418050c0603ed03090a00010405050903817d090a0001050e032e09160001060b0300090200010418050d0603d20209040001090e000001010405000902bab2010000000000039901010408050d0a03f30609060001040505000603f3770908000106039301090c00010421050903d602090200010405051403ea7c090400010427052d03ef03090800010405052303d17c090800010603ed7e090400010418050c0603ed03090a00010405050903817d090a0001050e032e09160001060b0300090200010418050d0603d20209040001090e0000010104090009022cb301000000000003cf110105090a03ec0109000001091600000101042200090242b301000000000003820101040905090a03f20a090a00010422051e038f75090200010409050903f10a09020001041f050503a376091000010409050903cf0d090c0001041f050c03fd7209140001050006039c7d09020001050c03e40209040001039c7d09020001042005090603a60a09020001041f051403c07809020001050006039a7d090a0001051403e60209020001040905090603910b09080001041f051403ef740906000104090509038f0909020001041f051503f2760914000104090509038e0909020001041f03f776091600010422050f03977e09040001060b0300090800010904000001010405000902e4b3010000000000039901010408050d0a03f30609060001040505000603f3770908000106039401090800010421050903d502090200010405051403ea7c090400010603ad7f09080001052306032a0902000103ea00090800010603ec7e090400010418050c0603ed03090a00010405050903817d090a0001050e032e09160001060b0300090200010418050d0603d20209040001090e00000101004743433a2028292031322e322e30004c696e6b65723a204c4c442031362e302e3200000000000000000000000000000000000000000000000000010000000400f1ff000000000000000000000000000000002200000000000400289a02000000000000000000000000002b00000002000300e23401000000000064000000000000000000000000000300e23401000000000000000000000000000000000000000300e43401000000000000000000000000000000000000000300ec340100000000000000000000000000fc00000000000300f83401000000000000000000000000000801000002000300f2b70100000000005600000000000000670100000200030002650100000000000800000000000000000000000000030046350100000000000000000000000000760100000200030046350100000000001000000000000000000000000000030046350100000000000000000000000000000000000000030056350100000000000000000000000000c7010000020003005635010000000000ee0000000000000000000000000003005635010000000000000000000000000000000000000003005835010000000000000000000000000000000000000003006235010000000000000000000000000042020000000003002e3601000000000000000000000000004e0200000100010072090100000000002b000000000000007802000002000300a4a90100000000000e00000000000000000000000000030044360100000000000000000000000000a5020000020003004436010000000000d404000000000000000000000000030044360100000000000000000000000000000000000000030046360100000000000000000000000000000000000000030060360100000000000000000000000000f8020000020003000245010000000000c600000000000000ce03000002000300f43b0100000000002c000000000000001f04000002000300203c0100000000002c000000000000007404000002000300183b010000000000dc000000000000008f05000000000300ae3a01000000000000000000000000009b05000001000100f90a0100000000003500000000000000c605000000000300bc3a0100000000000000000000000000d205000001000100d10a0100000000002800000000000000fd050000020003003ab20100000000000e000000000000006306000000000300d23a01000000000000000000000000006f06000000000300e83a01000000000000000000000000007b06000000000300f63a01000000000000000000000000008706000000000300003b01000000000000000000000000009306000001000100800a0100000000003000000000000000be060000000003000e3b01000000000000000000000000000000000000000300183b01000000000000000000000000000000000000000300183b010000000000000000000000000000000000000003001a3b01000000000000000000000000000000000000000300303b01000000000000000000000000000000000000000300f43b01000000000000000000000000000000000000000300f43b01000000000000000000000000000000000000000300f63b01000000000000000000000000000000000000000300f83b0100000000000000000000000000ca06000002000300fa640100000000000800000000000000d7060000020003001a650100000000000a000000000000000000000000000300203c01000000000000000000000000000000000000000300203c01000000000000000000000000000000000000000300223c01000000000000000000000000000000000000000300243c010000000000000000000000000000000000000003004c3c0100000000000000000000000000f2060000020003004c3c0100000000007a0100000000000000000000000003004c3c010000000000000000000000000000000000000003004e3c01000000000000000000000000000000000000000300663c010000000000000000000000000058070000000003008a3d01000000000000000000000000006407000001000100490b01000000000033000000000000008f07000000000300983d01000000000000000000000000009c070000010001007c0b0100000000002700000000000000c707000000000300a63d0100000000000000000000000000d407000000000300b03d0100000000000000000000000000e107000001000100a30b01000000000028000000000000000000000000000300c63d01000000000000000000000000000c08000002000300c63d010000000000aa010000000000000000000000000300c63d01000000000000000000000000000000000000000300c83d01000000000000000000000000000000000000000300e23d01000000000000000000000000007308000000000300383f01000000000000000000000000008008000001000100cb0b0100000000003200000000000000ab08000000000300463f0100000000000000000000000000b808000001000100fd0b0100000000002800000000000000e308000000000300503f0100000000000000000000000000f0080000000003005a3f01000000000000000000000000000000000000000300703f0100000000000000000000000000fd08000002000300703f010000000000c0010000000000000000000000000300703f01000000000000000000000000000000000000000300723f010000000000000000000000000000000000000003008c3f01000000000000000000000000006d090000000003000c4101000000000000000000000000007a09000001000100250c0100000000009100000000000000a5090000000003001a410100000000000000000000000000b209000001000100b60c0100000000002a00000000000000000000000000030030410100000000000000000000000000dd090000020003003041010000000000820100000000000000000000000003003041010000000000000000000000000000000000000003003241010000000000000000000000000000000000000003004c4101000000000000000000000000003b0a0000000003009c4201000000000000000000000000000000000000000300b2420100000000000000000000000000480a000002000300b24201000000000050020000000000000000000000000300b24201000000000000000000000000000000000000000300b44201000000000000000000000000000000000000000300ce420100000000000000000000000000960b000002000300d8c6010000000000680000000000000000000000000003000245010000000000000000000000000000000000000003000245010000000000000000000000000000000000000003000445010000000000000000000000000000000000000003001c4501000000000000000000000000000000000000000300c84501000000000000000000000000000000000000000300c84501000000000000000000000000000000000000000300cc4501000000000000000000000000000000000000000300004601000000000000000000000000000000000000000300004601000000000000000000000000000000000000000300024601000000000000000000000000005e0c000000000300024601000000000000000000000000006b0c000001000500789b0200000000001000000000000000940c000002000300eab50100000000004c00000000000000dc0c00000000030030470100000000000000000000000000e90c000001000100b7040100000000001100000000000000150d00000000030072470100000000000000000000000000220d0000000003009a4701000000000000000000000000002f0d000000000300dc470100000000000000000000000000390d0000000003002c480100000000000000000000000000460d0000000003006a480100000000000000000000000000530d00000000030090480100000000000000000000000000600d000002000300509a0100000000002200000000000000db0d000002000300f097010000000000d6000000000000006f0e000002000300729a0100000000003a00000000000000a80e000002000300a89b0100000000004200000000000000e70e0000000003002a490100000000000000000000000000f40e00000000030052490100000000000000000000000000010f000002000300ac9a010000000000fc00000000000000890f000002000300e4990100000000006c00000000000000bc0f000002000300ae9c01000000000064000000000000000f10000002000300a2a001000000000082000000000000005010000000000300ee4b01000000000000000000000000005d10000000000100600101000000000000000000000000006710000000000300fe4b01000000000000000000000000007110000002000300b23e0200000000005402000000000000a9100000020003003c6901000000000058000000000000000911000002000300e43a02000000000056020000000000004911000002000300ecba010000000000660100000000000090110000020003005e390200000000008601000000000000d111000000000300a84f0100000000000000000000000000db11000000000300ac4f0100000000000000000000000000e511000002000300426701000000000058000000000000003c12000002000300926601000000000058000000000000009812000002000300ea660100000000005800000000000000f212000002000300dc27020000000000ce020000000000002713000002000300e265010000000000580000000000000084130000020003003a660100000000005800000000000000df130000020003009a6701000000000058000000000000003a140000020003003265010000000000580000000000000095140000020003008a650100000000005800000000000000ee14000002000300229f01000000000072000000000000004415000002000300c8be010000000000b200000000000000c515000002000300f26701000000000052000000000000001e16000002000300dc2a02000000000018030000000000005516000002000300be6a0100000000004e00000000000000b616000002000300ec6901000000000086000000000000000217000002000300726a0100000000004c000000000000004e1700000200030094690100000000005800000000000000991700000200030044680100000000005800000000000000ec170000020003000c6b01000000000094000000000000004d180000020003006c4802000000000074000000000000007b18000002000300e048020000000000463a000000000000af1800000200030010350200000000004e04000000000000eb180000020003009c6801000000000052000000000000004b19000002000300f42d0200000000008c030000000000008f19000002000300ee680100000000004e00000000000000e219000002000300d2c0010000000000c0000000000000006e1a00000200030006410200000000006607000000000000ad1a00000200030080310200000000009003000000000000f41a0000020003003a3d0200000000007801000000000000291b000002000300a06b01000000000094000000000000008a1b00000000030074630100000000000000000000000000971b00000000030082630100000000000000000000000000a41b00000100010000020100000000001c00000000000000aa1b0000000003008c630100000000000000000000000000b51b000002000300a0a20100000000000e00000000000000e61b00000000030096630100000000000000000000000000f31b000001000100ee090100000000002b000000000000001e1c0000000003009e6301000000000000000000000000002b1c00000100010020020100000000002000000000000000551c000000000300ae630100000000000000000000000000621c000000000300b66301000000000000000000000000006f1c000001000100600201000000000020000000000000009a1c00000200030054ab0100000000000e00000000000000cd1c000000000300ce630100000000000000000000000000da1c000000000300d8630100000000000000000000000000e71c000000000300f2630100000000000000000000000000f41c000000000300fa630100000000000000000000000000011d000001000100400201000000000020000000000000002b1d0000000003000a640100000000000000000000000000381d00000000030012640100000000000000000000000000451d0000000003001c640100000000000000000000000000521d000000000300246401000000000000000000000000005f1d0000000003002e6401000000000000000000000000006c1d00000000030036640100000000000000000000000000791d00000000030040640100000000000000000000000000861d000001000100b00a010000000000210000000000000000000000000003004e640100000000000000000000000000b11d0000020003004e640100000000000a0000000000000000000000000003004e640100000000000000000000000000c31d00000200030084a20100000000001800000000000000000000000000030058640100000000000000000000000000f81d00000200030058640100000000000a00000000000000000000000000030058640100000000000000000000000000000000000000030062640100000000000000000000000000271e00000200030062640100000000000a0000000000000000000000000003006264010000000000000000000000000000000000000003006c640100000000000000000000000000301e0000020003006c64010000000000080000000000000000000000000003006c6401000000000000000000000000003b1e0000020003002a90010000000000d403000000000000000000000000030074640100000000000000000000000000c61e00000200030074640100000000000800000000000000000000000000030074640100000000000000000000000000d31e000002000300fe93010000000000f20300000000000000000000000003007c640100000000000000000000000000601f0000020003007c640100000000004e0000000000000000000000000003007c64010000000000000000000000000000000000000003007e6401000000000000000000000000000000000000000300886401000000000000000000000000000000000000000300ca6401000000000000000000000000006d1f000002000300ca6401000000000030000000000000000000000000000300ca6401000000000000000000000000000000000000000300cc6401000000000000000000000000000000000000000300d26401000000000000000000000000000000000000000300fa6401000000000000000000000000000000000000000300fa64010000000000000000000000000000000000000003000265010000000000000000000000000000000000000003000265010000000000000000000000000000000000000003000a6501000000000000000000000000007f1f0000020003000a65010000000000080000000000000000000000000003000a6501000000000000000000000000000000000000000300126501000000000000000000000000008e1f0000020003001265010000000000080000000000000000000000000003001265010000000000000000000000000000000000000003001a65010000000000000000000000000000000000000003001a650100000000000000000000000000000000000000030024650100000000000000000000000000a21f00000200030024650100000000000e00000000000000000000000000030024650100000000000000000000000000000000000000030024650100000000000000000000000000000000000000030024650100000000000000000000000000000000000000030026650100000000000000000000000000000000000000030026650100000000000000000000000000000000000000030028650100000000000000000000000000000000000000030032650100000000000000000000000000000000000000030032650100000000000000000000000000000000000000030032650100000000000000000000000000000000000000030034650100000000000000000000000000000000000000030038650100000000000000000000000000db1f000002000300acbd010000000000a20000000000000078200000000003006a65010000000000000000000000000085200000000003007265010000000000000000000000000000000000000003008a65010000000000000000000000000000000000000003008a65010000000000000000000000000000000000000003008c6501000000000000000000000000000000000000000300906501000000000000000000000000009220000000000300c26501000000000000000000000000009f20000000000300ca6501000000000000000000000000000000000000000300e26501000000000000000000000000000000000000000300e26501000000000000000000000000000000000000000300e46501000000000000000000000000000000000000000300e8650100000000000000000000000000ac200000000003001a660100000000000000000000000000b9200000000003002266010000000000000000000000000000000000000003003a66010000000000000000000000000000000000000003003a66010000000000000000000000000000000000000003003c660100000000000000000000000000000000000000030040660100000000000000000000000000c62000000000030072660100000000000000000000000000d3200000000003007a660100000000000000000000000000000000000000030092660100000000000000000000000000000000000000030092660100000000000000000000000000000000000000030094660100000000000000000000000000000000000000030098660100000000000000000000000000e020000000000300ca660100000000000000000000000000ed20000000000300d26601000000000000000000000000000000000000000300ea6601000000000000000000000000000000000000000300ea6601000000000000000000000000000000000000000300ec6601000000000000000000000000000000000000000300f0660100000000000000000000000000fa200000000003002267010000000000000000000000000007210000000003002a67010000000000000000000000000000000000000003004267010000000000000000000000000000000000000003004267010000000000000000000000000000000000000003004467010000000000000000000000000000000000000003004867010000000000000000000000000014210000000003007a67010000000000000000000000000021210000000003008267010000000000000000000000000000000000000003009a67010000000000000000000000000000000000000003009a67010000000000000000000000000000000000000003009c6701000000000000000000000000000000000000000300a06701000000000000000000000000002e21000000000300d26701000000000000000000000000003b21000000000300da6701000000000000000000000000000000000000000300f26701000000000000000000000000000000000000000300f26701000000000000000000000000000000000000000300f46701000000000000000000000000000000000000000300f667010000000000000000000000000048210000020003002ebd0100000000007e00000000000000cd2100000000030024680100000000000000000000000000da210000000003002c68010000000000000000000000000000000000000003004468010000000000000000000000000000000000000003004468010000000000000000000000000000000000000003004668010000000000000000000000000000000000000003004a680100000000000000000000000000e7210000000003007c680100000000000000000000000000f4210000000003008468010000000000000000000000000000000000000003009c68010000000000000000000000000000000000000003009c68010000000000000000000000000000000000000003009e6801000000000000000000000000000000000000000300a06801000000000000000000000000000122000002000300b6bc01000000000078000000000000008722000000000300ce6801000000000000000000000000009422000000000300d66801000000000000000000000000000000000000000300ee6801000000000000000000000000000000000000000300ee6801000000000000000000000000000000000000000300f06801000000000000000000000000000000000000000300f4680100000000000000000000000000a1220000000003001a690100000000000000000000000000ae220000000003002269010000000000000000000000000000000000000003003c69010000000000000000000000000000000000000003003c69010000000000000000000000000000000000000003003e690100000000000000000000000000000000000000030042690100000000000000000000000000bb2200000000030074690100000000000000000000000000c8220000000003007c69010000000000000000000000000000000000000003009469010000000000000000000000000000000000000003009469010000000000000000000000000000000000000003009669010000000000000000000000000000000000000003009a690100000000000000000000000000d522000000000300cc690100000000000000000000000000e222000000000300d46901000000000000000000000000000000000000000300ec6901000000000000000000000000000000000000000300ec6901000000000000000000000000000000000000000300ee6901000000000000000000000000000000000000000300f4690100000000000000000000000000ef22000002000300f2b901000000000062000000000000002823000002000300bcba01000000000030000000000000006823000000000300526a010000000000000000000000000075230000000003005c6a01000000000000000000000000000000000000000300726a01000000000000000000000000000000000000000300726a01000000000000000000000000000000000000000300746a01000000000000000000000000000000000000000300786a010000000000000000000000000082230000000003009c6a01000000000000000000000000008f23000000000300a46a01000000000000000000000000000000000000000300be6a01000000000000000000000000000000000000000300be6a01000000000000000000000000000000000000000300c06a01000000000000000000000000000000000000000300c46a01000000000000000000000000009c23000000000300ea6a0100000000000000000000000000a923000000000300f26a010000000000000000000000000000000000000003000c6b010000000000000000000000000000000000000003000c6b010000000000000000000000000000000000000003000e6b01000000000000000000000000000000000000000300126b0100000000000000000000000000b62300000200030052bc0100000000006400000000000000fb23000000000300686b01000000000000000000000000000824000000000300706b01000000000000000000000000001524000000000300806b01000000000000000000000000002224000000000300886b01000000000000000000000000000000000000000300a06b01000000000000000000000000000000000000000300a06b01000000000000000000000000000000000000000300a26b01000000000000000000000000000000000000000300a66b01000000000000000000000000002f24000000000300fc6b01000000000000000000000000003c24000000000300046c01000000000000000000000000004924000000000300146c010000000000000000000000000056240000000003001c6c01000000000000000000000000000000000000000300346c01000000000000000000000000006324000002000300346c010000000000bc000000000000000000000000000300346c01000000000000000000000000000000000000000300366c010000000000000000000000000000000000000003003e6c0100000000000000000000000000a624000002000300f06c0100000000009a00000000000000ec240000020003008a6d010000000000dc000000000000000000000000000300f06c01000000000000000000000000000000000000000300f06c01000000000000000000000000000000000000000300f26c01000000000000000000000000000000000000000300fa6c01000000000000000000000000002e25000000000300106d01000000000000000000000000003b25000001000100a002010000000000400000000000000000000000000003008a6d010000000000000000000000000000000000000003008a6d010000000000000000000000000000000000000003008e6d010000000000000000000000000000000000000003009a6d01000000000000000000000000007925000002000300666e010000000000ee1a0000000000000000000000000300666e0100000000000000000000000000bd25000000000400309a0200000000000000000000000000c725000000000400389a0200000000000000000000000000d125000000000400409a0200000000000000000000000000db25000000000400489a0200000000000000000000000000e525000000000400509a0200000000000000000000000000ef25000000000400589a0200000000000000000000000000f925000000000400609a02000000000000000000000000000326000000000400689a02000000000000000000000000000000000000000300666e01000000000000000000000000000000000000000300686e01000000000000000000000000000000000000000300826e01000000000000000000000000000d26000000000300026f01000000000000000000000000001a26000000000300166f01000000000000000000000000002726000000000300626f01000000000000000000000000003426000000000300766f01000000000000000000000000004126000000000300c06f01000000000000000000000000004e26000000000300da6f01000000000000000000000000005b260000000003002070010000000000000000000000000068260000000003003670010000000000000000000000000000000000000003005489010000000000000000000000000075260000020003005489010000000000f00000000000000000000000000003005489010000000000000000000000000000000000000003005689010000000000000000000000000000000000000003005e8901000000000000000000000000000000000000000300448a0100000000000000000000000000b326000002000300448a01000000000014040000000000000000000000000300448a01000000000000000000000000000000000000000300468a01000000000000000000000000000000000000000300608a0100000000000000000000000000f526000002000300588e0100000000003c000000000000002f27000000000300268b01000000000000000000000000003d27000001000100c0030100000000001c0000000000000046270000020003009e8e0100000000004c000000000000007f27000002000300ea8e0100000000004c00000000000000ca2700000200030062ab0100000000000e00000000000000fd270000000003009e8d01000000000000000000000000000b28000000000300b28d01000000000000000000000000001928000000000300bc8d01000000000000000000000000002728000000000300c68d01000000000000000000000000003428000000000300d08d01000000000000000000000000004228000001000100600301000000000021000000000000004b28000000000300da8d01000000000000000000000000005928000001000100900301000000000024000000000000006228000000000300e88d01000000000000000000000000007028000000000300f28d01000000000000000000000000007e28000001000100300301000000000021000000000000008728000000000300fc8d01000000000000000000000000009528000000000300068e0100000000000000000000000000a328000000000300108e0100000000000000000000000000b12800000100010000030100000000002300000000000000ba280000000003001e8e0100000000000000000000000000c72800000100010000040100000000001000000000000000f228000000000300388e01000000000000000000000000000029000001000100480401000000000010000000000000002b29000002000300948e0100000000000a0000000000000061290000000003004a8e01000000000000000000000000000000000000000300588e01000000000000000000000000000000000000000300588e01000000000000000000000000006f29000000000300708e01000000000000000000000000007d290000000003007e8e01000000000000000000000000000000000000000300948e01000000000000000000000000000000000000000300948e010000000000000000000000000000000000000003009e8e010000000000000000000000000000000000000003009e8e01000000000000000000000000008b29000000000300bc8e01000000000000000000000000009929000000000300c68e0100000000000000000000000000a729000000000300d48e01000000000000000000000000000000000000000300ea8e01000000000000000000000000000000000000000300ea8e0100000000000000000000000000b5290000000003000a8f0100000000000000000000000000c329000000000300148f0100000000000000000000000000d1290000000003002a8f0100000000000000000000000000df2900000100010058040100000000000d000000000000000000000000000300368f01000000000000000000000000000a2a000002000300368f010000000000f4000000000000000000000000000300368f0100000000000000000000000000492a00000000030002900100000000000000000000000000572a00000000030016900100000000000000000000000000652a0000000003002090010000000000000000000000000000000000000003002a90010000000000000000000000000000000000000003002a90010000000000000000000000000000000000000003002c900100000000000000000000000000000000000000030044900100000000000000000000000000732a0000000003004a900100000000000000000000000000812a000001000500d09a020000000000a800000000000000a92a00000000030056900100000000000000000000000000b72a00000000030000920100000000000000000000000000c52a00000000030042920100000000000000000000000000d32a00000000030072930100000000000000000000000000e12a0000000003007c930100000000000000000000000000ef2a0000000003008a930100000000000000000000000000fd2a0000000003009e9301000000000000000000000000000b2b000000000300a8930100000000000000000000000000192b000000000300bc930100000000000000000000000000272b000000000300c4930100000000000000000000000000352b000001000100e00201000000000020000000000000005f2b000000000300ce9301000000000000000000000000006d2b000000000300d69301000000000000000000000000007b2b000000000300e0930100000000000000000000000000892b000000000300e89301000000000000000000000000000000000000000300fe9301000000000000000000000000000000000000000300fe93010000000000000000000000000000000000000003000094010000000000000000000000000000000000000003001a940100000000000000000000000000972b0000000003001a940100000000000000000000000000a52b00000000030038940100000000000000000000000000b32b00000000030084940100000000000000000000000000c12b0000000003002c950100000000000000000000000000cf2b0000000003007c970100000000000000000000000000dd2b00000000030086970100000000000000000000000000eb2b00000000030094970100000000000000000000000000f92b000000000300a8970100000000000000000000000000072c000000000300c0970100000000000000000000000000152c000000000300c8970100000000000000000000000000232c000000000300d2970100000000000000000000000000312c000000000300da9701000000000000000000000000000000000000000300f09701000000000000000000000000000000000000000300f09701000000000000000000000000000000000000000300f29701000000000000000000000000000000000000000300009801000000000000000000000000003f2c000002000300c6980100000000004a00000000000000872c00000200030010990100000000003200000000000000e12c000000000300a4980100000000000000000000000000ef2c000001000100700401000000000019000000000000000000000000000300c69801000000000000000000000000000000000000000300c69801000000000000000000000000000000000000000300c89801000000000000000000000000000000000000000300cc980100000000000000000000000000000000000000030010990100000000000000000000000000000000000000030010990100000000000000000000000000000000000000030012990100000000000000000000000000000000000000030014990100000000000000000000000000f82c00000200030042990100000000006e0000000000000000000000000003004299010000000000000000000000000000000000000003004299010000000000000000000000000000000000000003004499010000000000000000000000000000000000000003004a990100000000000000000000000000432d00000200030022b501000000000062000000000000000000000000000300b0990100000000000000000000000000762d000002000300b09901000000000034000000000000000000000000000300b09901000000000000000000000000000000000000000300b29901000000000000000000000000000000000000000300b49901000000000000000000000000000000000000000300e49901000000000000000000000000000000000000000300e49901000000000000000000000000000000000000000300e69901000000000000000000000000000000000000000300f29901000000000000000000000000000000000000000300509a01000000000000000000000000000000000000000300509a01000000000000000000000000000000000000000300729a01000000000000000000000000000000000000000300729a01000000000000000000000000000000000000000300749a010000000000000000000000000000000000000003007a9a01000000000000000000000000000000000000000300ac9a01000000000000000000000000000000000000000300ac9a01000000000000000000000000000000000000000300ae9a01000000000000000000000000000000000000000300bc9a0100000000000000000000000000c32d000000000300d89a0100000000000000000000000000d12d000001000100ac040100000000000b00000000000000fd2d000000000300349b01000000000000000000000000000b2e0000000003008e9b01000000000000000000000000000000000000000300a89b01000000000000000000000000000000000000000300a89b01000000000000000000000000000000000000000300ea9b0100000000000000000000000000192e000002000300ea9b01000000000050000000000000000000000000000300ea9b01000000000000000000000000000000000000000300ec9b01000000000000000000000000000000000000000300f89b010000000000000000000000000000000000000003003a9c0100000000000000000000000000fc2e0000020003003a9c010000000000740000000000000000000000000003003a9c010000000000000000000000000000000000000003003c9c01000000000000000000000000000000000000000300449c0100000000000000000000000000d02f00000200030054b401000000000052000000000000007c300000000003009a9c01000000000000000000000000008a3000000100010090040100000000001c000000000000000000000000000300ae9c01000000000000000000000000000000000000000300ae9c01000000000000000000000000000000000000000300b09c01000000000000000000000000000000000000000300bc9c01000000000000000000000000000000000000000300129d01000000000000000000000000009330000002000300129d0100000000007a000000000000000000000000000300129d01000000000000000000000000000000000000000300149d010000000000000000000000000000000000000003001c9d010000000000000000000000000000000000000003008c9d01000000000000000000000000001b310000020003008c9d010000000000960100000000000000000000000003008c9d010000000000000000000000000000000000000003008e9d01000000000000000000000000000000000000000300a29d0100000000000000000000000000a531000000000300fa9e0100000000000000000000000000b331000000000300049f0100000000000000000000000000c1310000000003000e9f01000000000000000000000000000000000000000300229f01000000000000000000000000000000000000000300229f01000000000000000000000000000000000000000300949f0100000000000000000000000000cf31000002000300949f01000000000092000000000000000000000000000300949f01000000000000000000000000000000000000000300969f01000000000000000000000000000000000000000300989f01000000000000000000000000002a320000000003009c9f01000000000000000000000000003832000000000100880101000000000000000000000000004232000000000300aa9f01000000000000000000000000004b32000000000300b09f0100000000000000000000000000593200000100010043050100000000000f000000000000008432000000000300bc9f01000000000000000000000000008d32000000000300c29f01000000000000000000000000009b3200000100010038050100000000000b00000000000000c632000000000300ce9f0100000000000000000000000000cf32000000000300d29f0100000000000000000000000000dd3200000100010008050100000000000f000000000000000833000000000300da9f01000000000000000000000000001633000001000100180501000000000020000000000000004133000000000300e69f01000000000000000000000000004a33000000000300ec9f01000000000000000000000000005833000000000300fc9f0100000000000000000000000000613300000000030000a001000000000000000000000000006f33000001000100c80401000000000007000000000000009a3300000000030008a00100000000000000000000000000a833000001000100d0040100000000002000000000000000d333000002000300a2b10100000000009800000000000000000000000000030026a00100000000000000000000000000193400000200030026a00100000000000200000000000000000000000000030026a00100000000000000000000000000000000000000030028a00100000000000000000000000000583400000200030028a00100000000007a00000000000000000000000000030028a0010000000000000000000000000000000000000003002aa0010000000000000000000000000000000000000003002ea001000000000000000000000000000000000000000300a2a001000000000000000000000000000000000000000300a2a001000000000000000000000000000000000000000300a4a001000000000000000000000000000000000000000300a8a00100000000000000000000000000000000000000030024a10100000000000000000000000000993400000200030024a10100000000006001000000000000000000000000030024a10100000000000000000000000000000000000000030028a1010000000000000000000000000000000000000003004ca10100000000000000000000000000000000000000030084a20100000000000000000000000000000000000000030084a2010000000000000000000000000000000000000003009ca20100000000000000000000000000d5340000020003009ca2010000000000040000000000000000000000000003009ca2010000000000000000000000000000000000000003009ca2010000000000000000000000000000000000000003009ca2010000000000000000000000000000000000000003009ca2010000000000000000000000000000000000000003009ea2010000000000000000000000000000000000000003009ea201000000000000000000000000000000000000000300a0a201000000000000000000000000000000000000000300a0a201000000000000000000000000000000000000000300a0a201000000000000000000000000000000000000000300a0a201000000000000000000000000000000000000000300a0a201000000000000000000000000000000000000000300a0a201000000000000000000000000000000000000000300a2a201000000000000000000000000000000000000000300a2a201000000000000000000000000000000000000000300a4a201000000000000000000000000000000000000000300aea201000000000000000000000000000000000000000300aea201000000000000000000000000001035000002000300aea201000000000002000000000000000000000000000300aea201000000000000000000000000000000000000000300aea201000000000000000000000000000000000000000300aea201000000000000000000000000000000000000000300aea201000000000000000000000000000000000000000300b0a201000000000000000000000000000000000000000300b0a201000000000000000000000000009a35000000000400709a0200000000000000000000000000a435000002000300b0a201000000000042010000000000000000000000000300b0a201000000000000000000000000000000000000000300b0a201000000000000000000000000000000000000000300b0a201000000000000000000000000000000000000000300b2a201000000000000000000000000000000000000000300b4a201000000000000000000000000000000000000000300b6a20100000000000000000000000000d535000000000300c2a20100000000000000000000000000e335000001000100b805010000000000c8000000000000000000000000000300cea201000000000000000000000000000000000000000300d2a201000000000000000000000000000f36000000000300d6a201000000000000000000000000000000000000000300f6a201000000000000000000000000000000000000000300f8a20100000000000000000000000000000000000000030006a30100000000000000000000000000000000000000030020a30100000000000000000000000000000000000000030020a30100000000000000000000000000000000000000030022a30100000000000000000000000000000000000000030022a30100000000000000000000000000000000000000030026a30100000000000000000000000000000000000000030026a3010000000000000000000000000000000000000003002aa3010000000000000000000000000000000000000003002aa30100000000000000000000000000000000000000030032a30100000000000000000000000000000000000000030032a30100000000000000000000000000000000000000030034a30100000000000000000000000000000000000000030034a3010000000000000000000000000000000000000003003ca3010000000000000000000000000000000000000003003ca3010000000000000000000000000000000000000003003ea3010000000000000000000000000000000000000003003ea30100000000000000000000000000000000000000030042a30100000000000000000000000000000000000000030042a3010000000000000000000000000000000000000003004aa3010000000000000000000000000000000000000003004aa30100000000000000000000000000000000000000030050a30100000000000000000000000000000000000000030054a30100000000000000000000000000000000000000030058a30100000000000000000000000000000000000000030074a30100000000000000000000000000000000000000030078a3010000000000000000000000000000000000000003007aa3010000000000000000000000000000000000000003007aa3010000000000000000000000000000000000000003007ca3010000000000000000000000000000000000000003007ca30100000000000000000000000000000000000000030088a30100000000000000000000000000000000000000030088a3010000000000000000000000000000000000000003008aa3010000000000000000000000000000000000000003008aa30100000000000000000000000000000000000000030094a30100000000000000000000000000000000000000030094a30100000000000000000000000000000000000000030096a3010000000000000000000000000000000000000003009aa301000000000000000000000000000000000000000300a2a301000000000000000000000000000000000000000300a2a301000000000000000000000000000000000000000300a4a301000000000000000000000000000000000000000300a4a301000000000000000000000000000000000000000300aea301000000000000000000000000000000000000000300b0a301000000000000000000000000000000000000000300b4a301000000000000000000000000000000000000000300b4a301000000000000000000000000000000000000000300b6a301000000000000000000000000000000000000000300b6a301000000000000000000000000000000000000000300c2a301000000000000000000000000000000000000000300c2a301000000000000000000000000000000000000000300c4a301000000000000000000000000000000000000000300c4a301000000000000000000000000000000000000000300cca301000000000000000000000000000000000000000300cca301000000000000000000000000000000000000000300d0a301000000000000000000000000000000000000000300d0a301000000000000000000000000000000000000000300d6a301000000000000000000000000000000000000000300d6a301000000000000000000000000001d36000000000300d8a301000000000000000000000000002b36000001000100c00901000000000000000000000000000000000000000300d8a301000000000000000000000000005636000002000300f2a3010000000000e4010000000000000000000000000300eca301000000000000000000000000000000000000000300eea301000000000000000000000000000000000000000300f2a301000000000000000000000000000000000000000300f2a301000000000000000000000000000000000000000300f2a301000000000000000000000000000000000000000300f2a301000000000000000000000000000000000000000300f2a301000000000000000000000000000000000000000300f4a3010000000000000000000000000000000000000003000ea40100000000000000000000000000000000000000030010a40100000000000000000000000000000000000000030010a4010000000000000000000000000000000000000003001ca4010000000000000000000000000000000000000003001ca40100000000000000000000000000000000000000030028a4010000000000000000000000000000000000000003002ca4010000000000000000000000000000000000000003002ca40100000000000000000000000000000000000000030030a40100000000000000000000000000000000000000030030a40100000000000000000000000000000000000000030032a40100000000000000000000000000000000000000030034a40100000000000000000000000000000000000000030036a40100000000000000000000000000000000000000030038a4010000000000000000000000000000000000000003003ca4010000000000000000000000000000000000000003003ea4010000000000000000000000000000000000000003003ea40100000000000000000000000000000000000000030042a40100000000000000000000000000000000000000030042a40100000000000000000000000000000000000000030046a4010000000000000000000000000000000000000003004aa4010000000000000000000000000000000000000003004aa4010000000000000000000000000000000000000003004ca4010000000000000000000000000000000000000003004ca40100000000000000000000000000000000000000030054a40100000000000000000000000000000000000000030054a40100000000000000000000000000000000000000030056a40100000000000000000000000000000000000000030056a40100000000000000000000000000000000000000030058a40100000000000000000000000000000000000000030058a4010000000000000000000000000000000000000003005aa4010000000000000000000000000000000000000003005aa4010000000000000000000000000000000000000003005ca4010000000000000000000000000000000000000003005ea40100000000000000000000000000000000000000030060a40100000000000000000000000000000000000000030064a40100000000000000000000000000000000000000030068a40100000000000000000000000000000000000000030068a4010000000000000000000000000000000000000003006aa4010000000000000000000000000000000000000003006aa4010000000000000000000000000000000000000003006ca4010000000000000000000000000000000000000003006ca40100000000000000000000000000000000000000030072a40100000000000000000000000000000000000000030072a40100000000000000000000000000000000000000030076a40100000000000000000000000000000000000000030076a4010000000000000000000000000000000000000003007ca4010000000000000000000000000000000000000003007ca401000000000000000000000000008f36000002000300d6a5010000000000560000000000000000000000000003009ca401000000000000000000000000000000000000000300b8a401000000000000000000000000000000000000000300bca401000000000000000000000000000000000000000300e2a401000000000000000000000000000000000000000300e2a401000000000000000000000000000000000000000300e8a401000000000000000000000000000000000000000300e8a401000000000000000000000000000000000000000300eca401000000000000000000000000000000000000000300eca401000000000000000000000000000000000000000300f6a401000000000000000000000000000000000000000300f6a401000000000000000000000000000000000000000300faa401000000000000000000000000000000000000000300faa401000000000000000000000000000000000000000300fea401000000000000000000000000000000000000000300fea40100000000000000000000000000000000000000030012a50100000000000000000000000000000000000000030014a50100000000000000000000000000000000000000030014a5010000000000000000000000000000000000000003001aa5010000000000000000000000000000000000000003001aa5010000000000000000000000000000000000000003001ea5010000000000000000000000000000000000000003001ea5010000000000000000000000000000000000000003002ea5010000000000000000000000000000000000000003002ea50100000000000000000000000000000000000000030030a50100000000000000000000000000000000000000030030a50100000000000000000000000000000000000000030034a50100000000000000000000000000000000000000030038a5010000000000000000000000000000000000000003003aa50100000000000000000000000000000000000000030040a5010000000000000000000000000000000000000003004ca50100000000000000000000000000000000000000030050a50100000000000000000000000000000000000000030050a50100000000000000000000000000000000000000030052a50100000000000000000000000000000000000000030052a50100000000000000000000000000000000000000030054a50100000000000000000000000000000000000000030054a50100000000000000000000000000000000000000030060a50100000000000000000000000000000000000000030060a5010000000000000000000000000000000000000003006aa5010000000000000000000000000000000000000003006ea50100000000000000000000000000000000000000030082a50100000000000000000000000000000000000000030090a50100000000000000000000000000000000000000030090a50100000000000000000000000000000000000000030098a50100000000000000000000000000000000000000030098a501000000000000000000000000000000000000000300a0a501000000000000000000000000000000000000000300a0a501000000000000000000000000000000000000000300b0a501000000000000000000000000000000000000000300b0a501000000000000000000000000000000000000000300c0a501000000000000000000000000000000000000000300c2a501000000000000000000000000000000000000000300c6a501000000000000000000000000000000000000000300cea501000000000000000000000000000000000000000300d0a501000000000000000000000000000000000000000300d0a501000000000000000000000000000000000000000300d6a501000000000000000000000000000000000000000300d6a501000000000000000000000000000000000000000300d6a501000000000000000000000000000000000000000300d6a501000000000000000000000000000000000000000300d6a501000000000000000000000000000000000000000300d6a501000000000000000000000000000000000000000300d8a501000000000000000000000000000000000000000300e2a501000000000000000000000000000000000000000300f2a501000000000000000000000000000000000000000300f6a50100000000000000000000000000000000000000030004a60100000000000000000000000000000000000000030006a60100000000000000000000000000000000000000030018a6010000000000000000000000000000000000000003001ca6010000000000000000000000000000000000000003001ea60100000000000000000000000000000000000000030028a6010000000000000000000000000000000000000003002ca6010000000000000000000000000000000000000003002ca60100000000000000000000000000d636000000000400789a0200000000000000000000000000e036000000000400809a0200000000000000000000000000ea360000020003002ca6010000000000780300000000000000000000000003002ca6010000000000000000000000000000000000000003002ca6010000000000000000000000000000000000000003002ca6010000000000000000000000000000000000000003002ea6010000000000000000000000000000000000000003002ea6010000000000000000000000000000000000000003002ea60100000000000000000000000000000000000000030040a60100000000000000000000000000000000000000030044a60100000000000000000000000000000000000000030044a60100000000000000000000000000000000000000030046a60100000000000000000000000000000000000000030046a6010000000000000000000000000000000000000003004ea6010000000000000000000000000000000000000003004ea60100000000000000000000000000000000000000030052a60100000000000000000000000000000000000000030056a6010000000000000000000000000000000000000003005aa6010000000000000000000000000000000000000003005aa6010000000000000000000000000000000000000003005ea6010000000000000000000000000000000000000003005ea60100000000000000000000000000000000000000030070a60100000000000000000000000000000000000000030070a60100000000000000000000000000000000000000030074a60100000000000000000000000000000000000000030074a60100000000000000000000000000000000000000030076a6010000000000000000000000000000000000000003007aa6010000000000000000000000000000000000000003007aa6010000000000000000000000000000000000000003007ea6010000000000000000000000000000000000000003007ea60100000000000000000000000000000000000000030080a60100000000000000000000000000000000000000030080a60100000000000000000000000000000000000000030082a60100000000000000000000000000000000000000030082a60100000000000000000000000000000000000000030086a60100000000000000000000000000000000000000030086a6010000000000000000000000000000000000000003008ea60100000000000000000000000000000000000000030092a60100000000000000000000000000000000000000030096a60100000000000000000000000000000000000000030096a6010000000000000000000000000000000000000003009aa6010000000000000000000000000000000000000003009aa6010000000000000000000000000000000000000003009ea6010000000000000000000000000000000000000003009ea601000000000000000000000000000000000000000300a2a601000000000000000000000000000000000000000300a6a601000000000000000000000000000000000000000300a6a601000000000000000000000000000000000000000300a8a601000000000000000000000000000000000000000300aca601000000000000000000000000000000000000000300b0a601000000000000000000000000000000000000000300b0a601000000000000000000000000000000000000000300b4a601000000000000000000000000000000000000000300b8a601000000000000000000000000000000000000000300bca601000000000000000000000000000000000000000300bca601000000000000000000000000000000000000000300bea601000000000000000000000000000000000000000300c2a601000000000000000000000000000000000000000300c6a601000000000000000000000000000000000000000300c6a601000000000000000000000000000000000000000300c8a601000000000000000000000000000000000000000300c8a601000000000000000000000000000000000000000300cca601000000000000000000000000000000000000000300cca601000000000000000000000000000000000000000300eaa601000000000000000000000000000000000000000300eaa601000000000000000000000000000000000000000300eea601000000000000000000000000000000000000000300eea601000000000000000000000000000000000000000300f2a601000000000000000000000000000000000000000300f6a601000000000000000000000000000000000000000300fea60100000000000000000000000000000000000000030002a70100000000000000000000000000000000000000030006a7010000000000000000000000000000000000000003000aa7010000000000000000000000000000000000000003000ea70100000000000000000000000000000000000000030012a70100000000000000000000000000000000000000030012a70100000000000000000000000000000000000000030016a70100000000000000000000000000000000000000030016a7010000000000000000000000000000000000000003001aa7010000000000000000000000000000000000000003001aa7010000000000000000000000000000000000000003001ea70100000000000000000000000000000000000000030022a70100000000000000000000000000000000000000030022a70100000000000000000000000000000000000000030028a7010000000000000000000000000000000000000003002ca7010000000000000000000000000000000000000003002ea7010000000000000000000000000000000000000003002ea70100000000000000000000000000000000000000030034a70100000000000000000000000000000000000000030034a70100000000000000000000000000000000000000030038a70100000000000000000000000000000000000000030038a7010000000000000000000000000000000000000003003aa7010000000000000000000000000000000000000003003ea7010000000000000000000000000000000000000003003ea70100000000000000000000000000000000000000030042a70100000000000000000000000000000000000000030042a7010000000000000000000000000000000000000003004aa7010000000000000000000000000000000000000003004aa7010000000000000000000000000000000000000003004ea7010000000000000000000000000000000000000003004ea70100000000000000000000000000000000000000030050a70100000000000000000000000000000000000000030050a70100000000000000000000000000000000000000030054a70100000000000000000000000000000000000000030054a70100000000000000000000000000000000000000030058a70100000000000000000000000000000000000000030058a7010000000000000000000000000000000000000003005aa7010000000000000000000000000000000000000003005aa7010000000000000000000000000000000000000003005ca7010000000000000000000000000000000000000003005ca70100000000000000000000000000000000000000030060a70100000000000000000000000000000000000000030064a7010000000000000000000000000000000000000003006ca7010000000000000000000000000000000000000003006ca70100000000000000000000000000000000000000030070a70100000000000000000000000000000000000000030072a70100000000000000000000000000000000000000030072a70100000000000000000000000000000000000000030076a70100000000000000000000000000000000000000030076a7010000000000000000000000000000000000000003007aa7010000000000000000000000000000000000000003007ea7010000000000000000000000000000000000000003007ea70100000000000000000000000000000000000000030080a70100000000000000000000000000000000000000030080a70100000000000000000000000000000000000000030088a70100000000000000000000000000000000000000030088a7010000000000000000000000000000000000000003008aa7010000000000000000000000000000000000000003008aa7010000000000000000000000000000000000000003008ca7010000000000000000000000000000000000000003008ca70100000000000000000000000000000000000000030090a70100000000000000000000000000000000000000030090a70100000000000000000000000000000000000000030096a70100000000000000000000000000000000000000030096a7010000000000000000000000000000000000000003009ea7010000000000000000000000000000000000000003009ea701000000000000000000000000000000000000000300a4a701000000000000000000000000000000000000000300a4a701000000000000000000000000000000000000000300a8a701000000000000000000000000000000000000000300a8a701000000000000000000000000000000000000000300aaa701000000000000000000000000000000000000000300aea701000000000000000000000000000000000000000300aea701000000000000000000000000000000000000000300b0a701000000000000000000000000000000000000000300b0a701000000000000000000000000000000000000000300b8a701000000000000000000000000000000000000000300b8a701000000000000000000000000000000000000000300baa701000000000000000000000000000000000000000300baa701000000000000000000000000000000000000000300bca701000000000000000000000000000000000000000300bca701000000000000000000000000000000000000000300bea701000000000000000000000000000000000000000300bea701000000000000000000000000000000000000000300c0a701000000000000000000000000000000000000000300c0a701000000000000000000000000000000000000000300c2a701000000000000000000000000000000000000000300c2a701000000000000000000000000000000000000000300c8a701000000000000000000000000000000000000000300cca701000000000000000000000000000000000000000300cca701000000000000000000000000000000000000000300cea701000000000000000000000000000000000000000300cea701000000000000000000000000000000000000000300d6a701000000000000000000000000000000000000000300d6a701000000000000000000000000000000000000000300d8a701000000000000000000000000000000000000000300d8a701000000000000000000000000000000000000000300daa701000000000000000000000000000000000000000300daa701000000000000000000000000000000000000000300dca701000000000000000000000000000000000000000300dca701000000000000000000000000001937000000000300e0a701000000000000000000000000002737000000000300e8a701000000000000000000000000000000000000000300fea70100000000000000000000000000000000000000030004a80100000000000000000000000000000000000000030012a80100000000000000000000000000000000000000030012a80100000000000000000000000000000000000000030016a80100000000000000000000000000000000000000030018a8010000000000000000000000000000000000000003001ca8010000000000000000000000000000000000000003001ea8010000000000000000000000000000000000000003001ea80100000000000000000000000000000000000000030022a80100000000000000000000000000000000000000030022a80100000000000000000000000000000000000000030024a80100000000000000000000000000000000000000030024a80100000000000000000000000000000000000000030026a80100000000000000000000000000000000000000030028a80100000000000000000000000000000000000000030028a8010000000000000000000000000000000000000003002aa80100000000000000000000000000000000000000030034a80100000000000000000000000000000000000000030038a8010000000000000000000000000000000000000003003ca8010000000000000000000000000000000000000003003ca80100000000000000000000000000000000000000030040a80100000000000000000000000000000000000000030040a80100000000000000000000000000000000000000030046a80100000000000000000000000000000000000000030046a80100000000000000000000000000000000000000030048a80100000000000000000000000000000000000000030048a8010000000000000000000000000000000000000003004ca8010000000000000000000000000000000000000003004ea80100000000000000000000000000000000000000030050a80100000000000000000000000000000000000000030050a80100000000000000000000000000000000000000030054a80100000000000000000000000000000000000000030056a80100000000000000000000000000000000000000030058a80100000000000000000000000000000000000000030058a8010000000000000000000000000000000000000003005aa8010000000000000000000000000000000000000003005aa8010000000000000000000000000000000000000003005ea8010000000000000000000000000000000000000003005ea80100000000000000000000000000000000000000030060a80100000000000000000000000000000000000000030060a80100000000000000000000000000000000000000030064a80100000000000000000000000000000000000000030066a80100000000000000000000000000000000000000030066a80100000000000000000000000000000000000000030068a80100000000000000000000000000000000000000030068a8010000000000000000000000000000000000000003006aa8010000000000000000000000000000000000000003006ea80100000000000000000000000000000000000000030072a80100000000000000000000000000000000000000030074a80100000000000000000000000000000000000000030076a80100000000000000000000000000000000000000030078a80100000000000000000000000000000000000000030078a8010000000000000000000000000000000000000003007aa8010000000000000000000000000000000000000003007aa8010000000000000000000000000000000000000003007ca8010000000000000000000000000000000000000003007ca80100000000000000000000000000000000000000030080a80100000000000000000000000000000000000000030080a80100000000000000000000000000000000000000030084a80100000000000000000000000000000000000000030086a80100000000000000000000000000000000000000030088a8010000000000000000000000000000000000000003008ca8010000000000000000000000000000000000000003008ca80100000000000000000000000000000000000000030090a80100000000000000000000000000000000000000030090a80100000000000000000000000000000000000000030092a80100000000000000000000000000000000000000030092a80100000000000000000000000000000000000000030098a80100000000000000000000000000000000000000030098a8010000000000000000000000000000000000000003009ca801000000000000000000000000000000000000000300a0a801000000000000000000000000000000000000000300a4a801000000000000000000000000000000000000000300aaa801000000000000000000000000000000000000000300b0a801000000000000000000000000000000000000000300b0a801000000000000000000000000000000000000000300b2a801000000000000000000000000000000000000000300b2a801000000000000000000000000000000000000000300b4a801000000000000000000000000000000000000000300b4a801000000000000000000000000000000000000000300b8a801000000000000000000000000000000000000000300baa801000000000000000000000000000000000000000300bca801000000000000000000000000000000000000000300c0a801000000000000000000000000000000000000000300c0a801000000000000000000000000000000000000000300c2a801000000000000000000000000000000000000000300c2a801000000000000000000000000000000000000000300c4a801000000000000000000000000000000000000000300c4a801000000000000000000000000000000000000000300c8a801000000000000000000000000000000000000000300c8a801000000000000000000000000000000000000000300caa801000000000000000000000000000000000000000300caa801000000000000000000000000000000000000000300cea801000000000000000000000000000000000000000300d0a801000000000000000000000000000000000000000300d4a801000000000000000000000000000000000000000300d6a801000000000000000000000000000000000000000300d6a801000000000000000000000000000000000000000300daa801000000000000000000000000000000000000000300daa801000000000000000000000000000000000000000300dca801000000000000000000000000000000000000000300dca801000000000000000000000000000000000000000300dea801000000000000000000000000000000000000000300dea801000000000000000000000000000000000000000300e2a801000000000000000000000000000000000000000300e2a801000000000000000000000000000000000000000300e8a801000000000000000000000000000000000000000300e8a801000000000000000000000000000000000000000300eca801000000000000000000000000000000000000000300eca801000000000000000000000000000000000000000300f2a801000000000000000000000000000000000000000300f2a80100000000000000000000000000000000000000030018a90100000000000000000000000000000000000000030018a9010000000000000000000000000000000000000003001ca90100000000000000000000000000000000000000030020a90100000000000000000000000000000000000000030022a90100000000000000000000000000000000000000030028a90100000000000000000000000000000000000000030036a9010000000000000000000000000000000000000003003aa9010000000000000000000000000000000000000003003aa9010000000000000000000000000000000000000003003ca9010000000000000000000000000000000000000003003ca9010000000000000000000000000000000000000003003ea9010000000000000000000000000000000000000003003ea9010000000000000000000000000000000000000003004aa9010000000000000000000000000000000000000003004aa90100000000000000000000000000000000000000030054a90100000000000000000000000000000000000000030058a90100000000000000000000000000000000000000030066a90100000000000000000000000000000000000000030066a9010000000000000000000000000000000000000003006ea9010000000000000000000000000000000000000003006ea90100000000000000000000000000000000000000030072a90100000000000000000000000000000000000000030072a90100000000000000000000000000000000000000030076a90100000000000000000000000000000000000000030076a90100000000000000000000000000000000000000030086a90100000000000000000000000000000000000000030088a90100000000000000000000000000000000000000030088a9010000000000000000000000000000000000000003008ca9010000000000000000000000000000000000000003008ca901000000000000000000000000000000000000000300a0a901000000000000000000000000000000000000000300a4a901000000000000000000000000000000000000000300a4a901000000000000000000000000000000000000000300a4a901000000000000000000000000000000000000000300a4a901000000000000000000000000000000000000000300a4a901000000000000000000000000000000000000000300a6a901000000000000000000000000000000000000000300a6a901000000000000000000000000000000000000000300a8a901000000000000000000000000000000000000000300b2a901000000000000000000000000000000000000000300b2a901000000000000000000000000003537000002000300b2a90100000000007e010000000000000000000000000300b2a901000000000000000000000000000000000000000300b2a901000000000000000000000000000000000000000300b2a901000000000000000000000000000000000000000300b4a901000000000000000000000000000000000000000300c4a901000000000000000000000000000000000000000300caa901000000000000000000000000000000000000000300caa901000000000000000000000000000000000000000300d2a901000000000000000000000000000000000000000300d2a901000000000000000000000000000000000000000300d6a901000000000000000000000000000000000000000300d6a901000000000000000000000000000000000000000300dea901000000000000000000000000000000000000000300dea901000000000000000000000000000000000000000300e0a901000000000000000000000000000000000000000300e4a901000000000000000000000000000000000000000300e4a901000000000000000000000000000000000000000300e8a901000000000000000000000000000000000000000300eca901000000000000000000000000005c3700000000030006aa010000000000000000000000000000000000000003000eaa010000000000000000000000000000000000000003000eaa0100000000000000000000000000000000000000030010aa0100000000000000000000000000000000000000030012aa0100000000000000000000000000000000000000030016aa010000000000000000000000000000000000000003001aaa0100000000000000000000000000000000000000030020aa0100000000000000000000000000000000000000030020aa0100000000000000000000000000000000000000030022aa0100000000000000000000000000000000000000030024aa0100000000000000000000000000000000000000030028aa010000000000000000000000000000000000000003002caa010000000000000000000000000000000000000003002eaa010000000000000000000000000000000000000003002eaa0100000000000000000000000000000000000000030032aa0100000000000000000000000000000000000000030032aa0100000000000000000000000000000000000000030034aa010000000000000000000000000000000000000003003aaa010000000000000000000000000000000000000003003aaa0100000000000000000000000000000000000000030040aa0100000000000000000000000000000000000000030040aa010000000000000000000000000000000000000003004aaa010000000000000000000000000000000000000003004eaa0100000000000000000000000000000000000000030050aa0100000000000000000000000000000000000000030052aa0100000000000000000000000000000000000000030052aa0100000000000000000000000000000000000000030054aa0100000000000000000000000000000000000000030058aa0100000000000000000000000000000000000000030060aa0100000000000000000000000000000000000000030060aa0100000000000000000000000000000000000000030066aa0100000000000000000000000000000000000000030066aa0100000000000000000000000000000000000000030070aa0100000000000000000000000000000000000000030074aa0100000000000000000000000000000000000000030076aa0100000000000000000000000000000000000000030078aa0100000000000000000000000000000000000000030078aa010000000000000000000000000000000000000003007aaa010000000000000000000000000000000000000003007eaa0100000000000000000000000000000000000000030080aa0100000000000000000000000000000000000000030080aa0100000000000000000000000000000000000000030084aa0100000000000000000000000000000000000000030084aa0100000000000000000000000000000000000000030086aa0100000000000000000000000000000000000000030088aa010000000000000000000000000000000000000003008caa010000000000000000000000000000000000000003008caa010000000000000000000000000000000000000003008eaa010000000000000000000000000000000000000003008eaa010000000000000000000000000000000000000003009eaa010000000000000000000000000000000000000003009eaa01000000000000000000000000000000000000000300a2aa01000000000000000000000000000000000000000300a2aa01000000000000000000000000000000000000000300a6aa01000000000000000000000000000000000000000300aeaa01000000000000000000000000000000000000000300c0aa01000000000000000000000000000000000000000300c0aa01000000000000000000000000000000000000000300c2aa01000000000000000000000000000000000000000300c4aa01000000000000000000000000000000000000000300c8aa01000000000000000000000000000000000000000300ccaa01000000000000000000000000000000000000000300d2aa01000000000000000000000000000000000000000300d2aa01000000000000000000000000000000000000000300d4aa01000000000000000000000000000000000000000300d8aa01000000000000000000000000000000000000000300dcaa01000000000000000000000000000000000000000300dcaa01000000000000000000000000000000000000000300deaa01000000000000000000000000000000000000000300deaa01000000000000000000000000000000000000000300e8aa01000000000000000000000000000000000000000300e8aa01000000000000000000000000000000000000000300ecaa01000000000000000000000000000000000000000300ecaa01000000000000000000000000000000000000000300f2aa01000000000000000000000000000000000000000300f2aa01000000000000000000000000000000000000000300f4aa01000000000000000000000000000000000000000300f8aa01000000000000000000000000000000000000000300f8aa01000000000000000000000000000000000000000300fcaa01000000000000000000000000000000000000000300fcaa0100000000000000000000000000000000000000030000ab0100000000000000000000000000000000000000030000ab0100000000000000000000000000000000000000030004ab0100000000000000000000000000000000000000030004ab0100000000000000000000000000000000000000030008ab0100000000000000000000000000000000000000030010ab0100000000000000000000000000000000000000030016ab010000000000000000000000000000000000000003001cab010000000000000000000000000000000000000003002cab0100000000000000000000000000000000000000030030ab0100000000000000000000000000000000000000030030ab01000000000000000000000000006a3700000200030030ab0100000000001200000000000000000000000000030030ab0100000000000000000000000000000000000000030030ab0100000000000000000000000000000000000000030030ab0100000000000000000000000000000000000000030030ab0100000000000000000000000000c43700000000030036ab0100000000000000000000000000d23700000100010053050100000000000b00000000000000000000000000030042ab0100000000000000000000000000000000000000030042ab0100000000000000000000000000000000000000030042ab0100000000000000000000000000fe3700000200030042ab0100000000001200000000000000000000000000030042ab0100000000000000000000000000000000000000030042ab0100000000000000000000000000000000000000030042ab0100000000000000000000000000000000000000030042ab01000000000000000000000000005b3800000000030048ab010000000000000000000000000069380000010001005e050100000000000e00000000000000000000000000030054ab0100000000000000000000000000000000000000030054ab0100000000000000000000000000000000000000030054ab0100000000000000000000000000000000000000030054ab0100000000000000000000000000000000000000030054ab0100000000000000000000000000000000000000030054ab0100000000000000000000000000000000000000030056ab0100000000000000000000000000000000000000030056ab0100000000000000000000000000000000000000030058ab0100000000000000000000000000000000000000030062ab0100000000000000000000000000000000000000030062ab0100000000000000000000000000000000000000030062ab0100000000000000000000000000000000000000030062ab0100000000000000000000000000000000000000030062ab0100000000000000000000000000000000000000030064ab0100000000000000000000000000000000000000030064ab0100000000000000000000000000000000000000030064ab0100000000000000000000000000000000000000030066ab0100000000000000000000000000000000000000030070ab0100000000000000000000000000000000000000030070ab0100000000000000000000000000000000000000030070ab0100000000000000000000000000953800000200030070ab0100000000007000000000000000000000000000030070ab0100000000000000000000000000000000000000030070ab0100000000000000000000000000000000000000030070ab0100000000000000000000000000000000000000030072ab0100000000000000000000000000000000000000030074ab0100000000000000000000000000000000000000030076ab0100000000000000000000000000000000000000030076ab010000000000000000000000000000000000000003007eab010000000000000000000000000000000000000003007eab0100000000000000000000000000000000000000030086ab0100000000000000000000000000000000000000030086ab0100000000000000000000000000000000000000030088ab0100000000000000000000000000000000000000030088ab010000000000000000000000000000000000000003008cab010000000000000000000000000000000000000003008cab0100000000000000000000000000000000000000030094ab0100000000000000000000000000000000000000030096ab0100000000000000000000000000000000000000030096ab010000000000000000000000000000000000000003009eab010000000000000000000000000000000000000003009eab01000000000000000000000000000000000000000300a2ab01000000000000000000000000000000000000000300a2ab01000000000000000000000000000000000000000300acab01000000000000000000000000000000000000000300acab01000000000000000000000000000000000000000300b6ab0100000000000000000000000000f538000000000300b6ab01000000000000000000000000000339000001000100b60501000000000002000000000000000000000000000300b6ab01000000000000000000000000000000000000000300ccab01000000000000000000000000000000000000000300ccab01000000000000000000000000000000000000000300ceab01000000000000000000000000000000000000000300d2ab01000000000000000000000000000000000000000300d2ab01000000000000000000000000000000000000000300e0ab01000000000000000000000000000000000000000300e0ab01000000000000000000000000000000000000000300e0ab01000000000000000000000000002f39000000000400889a02000000000000000000000000003939000000000400909a02000000000000000000000000004339000000000400989a02000000000000000000000000004d39000002000300e0ab010000000000bc010000000000000000000000000300e0ab01000000000000000000000000000000000000000300e0ab01000000000000000000000000000000000000000300e0ab01000000000000000000000000000000000000000300e2ab01000000000000000000000000000000000000000300fcab0100000000000000000000000000b53900000000030006ac0100000000000000000000000000c3390000000003000eac0100000000000000000000000000d13900000000030016ac0100000000000000000000000000000000000000030026ac0100000000000000000000000000000000000000030026ac0100000000000000000000000000df390000000003002eac010000000000000000000000000000000000000003003eac010000000000000000000000000000000000000003003eac0100000000000000000000000000000000000000030042ac0100000000000000000000000000000000000000030042ac010000000000000000000000000000000000000003004cac010000000000000000000000000000000000000003004cac0100000000000000000000000000000000000000030050ac010000000000000000000000000000000000000003005eac010000000000000000000000000000000000000003005eac0100000000000000000000000000000000000000030066ac0100000000000000000000000000000000000000030066ac0100000000000000000000000000000000000000030070ac0100000000000000000000000000000000000000030070ac0100000000000000000000000000000000000000030078ac0100000000000000000000000000000000000000030078ac010000000000000000000000000000000000000003007eac010000000000000000000000000000000000000003007eac0100000000000000000000000000000000000000030082ac0100000000000000000000000000000000000000030084ac0100000000000000000000000000000000000000030090ac0100000000000000000000000000000000000000030092ac0100000000000000000000000000000000000000030098ac0100000000000000000000000000000000000000030098ac01000000000000000000000000000000000000000300a0ac01000000000000000000000000000000000000000300a4ac01000000000000000000000000000000000000000300a4ac01000000000000000000000000000000000000000300b2ac01000000000000000000000000000000000000000300b8ac01000000000000000000000000000000000000000300bcac01000000000000000000000000000000000000000300bcac01000000000000000000000000000000000000000300c0ac01000000000000000000000000000000000000000300c0ac01000000000000000000000000000000000000000300c6ac01000000000000000000000000000000000000000300c8ac01000000000000000000000000000000000000000300c8ac01000000000000000000000000000000000000000300caac01000000000000000000000000000000000000000300caac01000000000000000000000000000000000000000300d2ac01000000000000000000000000000000000000000300d2ac01000000000000000000000000000000000000000300dcac01000000000000000000000000000000000000000300deac01000000000000000000000000000000000000000300deac01000000000000000000000000000000000000000300e0ac01000000000000000000000000000000000000000300e0ac01000000000000000000000000000000000000000300e8ac01000000000000000000000000000000000000000300e8ac01000000000000000000000000000000000000000300eaac01000000000000000000000000000000000000000300f0ac01000000000000000000000000000000000000000300f0ac01000000000000000000000000000000000000000300fcac01000000000000000000000000000000000000000300feac0100000000000000000000000000000000000000030002ad0100000000000000000000000000000000000000030002ad0100000000000000000000000000000000000000030006ad010000000000000000000000000000000000000003000aad0100000000000000000000000000000000000000030010ad0100000000000000000000000000000000000000030010ad010000000000000000000000000000000000000003001cad0100000000000000000000000000000000000000030024ad0100000000000000000000000000000000000000030024ad0100000000000000000000000000000000000000030026ad0100000000000000000000000000000000000000030028ad0100000000000000000000000000000000000000030030ad0100000000000000000000000000000000000000030030ad0100000000000000000000000000000000000000030032ad0100000000000000000000000000000000000000030032ad0100000000000000000000000000000000000000030036ad0100000000000000000000000000000000000000030036ad010000000000000000000000000000000000000003003aad010000000000000000000000000000000000000003003aad010000000000000000000000000000000000000003004ead0100000000000000000000000000000000000000030054ad0100000000000000000000000000000000000000030062ad010000000000000000000000000000000000000003006aad010000000000000000000000000000000000000003006aad010000000000000000000000000000000000000003006ead010000000000000000000000000000000000000003006ead010000000000000000000000000000000000000003007ead0100000000000000000000000000000000000000030098ad010000000000000000000000000000000000000003009cad010000000000000000000000000000000000000003009cad0100000000000000000000000000ed390000020003009cad010000000000b40000000000000000000000000003009cad010000000000000000000000000000000000000003009cad010000000000000000000000000000000000000003009cad010000000000000000000000000000000000000003009ead01000000000000000000000000000000000000000300a0ad01000000000000000000000000000000000000000300a8ad01000000000000000000000000000000000000000300aaad01000000000000000000000000000000000000000300aaad01000000000000000000000000000000000000000300aead01000000000000000000000000000000000000000300aead01000000000000000000000000000000000000000300b6ad01000000000000000000000000000000000000000300b6ad01000000000000000000000000000000000000000300bcad01000000000000000000000000000000000000000300bcad01000000000000000000000000000000000000000300c0ad01000000000000000000000000000000000000000300c8ad01000000000000000000000000000000000000000300ccad01000000000000000000000000000000000000000300d8ad01000000000000000000000000000000000000000300d8ad01000000000000000000000000000000000000000300dead01000000000000000000000000000000000000000300dead01000000000000000000000000000000000000000300e2ad01000000000000000000000000000000000000000300eaad01000000000000000000000000000000000000000300f0ad01000000000000000000000000000000000000000300f8ad01000000000000000000000000000000000000000300fcad0100000000000000000000000000000000000000030008ae010000000000000000000000000000000000000003000eae0100000000000000000000000000000000000000030016ae010000000000000000000000000000000000000003001cae0100000000000000000000000000000000000000030024ae010000000000000000000000000000000000000003002aae0100000000000000000000000000000000000000030032ae0100000000000000000000000000000000000000030036ae0100000000000000000000000000000000000000030040ae0100000000000000000000000000000000000000030040ae010000000000000000000000000000000000000003004aae010000000000000000000000000000000000000003004cae0100000000000000000000000000000000000000030050ae0100000000000000000000000000000000000000030050ae0100000000000000000000000000203a00000200030050ae0100000000003800000000000000000000000000030050ae0100000000000000000000000000000000000000030050ae0100000000000000000000000000000000000000030050ae0100000000000000000000000000000000000000030052ae0100000000000000000000000000000000000000030052ae0100000000000000000000000000000000000000030054ae0100000000000000000000000000513a0000000003006eae01000000000000000000000000005f3a00000100010080060100000000003000000000000000000000000000030082ae0100000000000000000000000000000000000000030084ae0100000000000000000000000000000000000000030088ae0100000000000000000000000000000000000000030088ae01000000000000000000000000008b3a00000200030088ae0100000000000a00000000000000000000000000030088ae0100000000000000000000000000000000000000030088ae0100000000000000000000000000000000000000030088ae0100000000000000000000000000000000000000030088ae0100000000000000000000000000000000000000030092ae0100000000000000000000000000000000000000030092ae0100000000000000000000000000e13a00000200030092ae010000000000b600000000000000000000000000030092ae0100000000000000000000000000000000000000030092ae0100000000000000000000000000000000000000030092ae0100000000000000000000000000000000000000030094ae0100000000000000000000000000000000000000030094ae0100000000000000000000000000000000000000030096ae01000000000000000000000000000000000000000300a0ae01000000000000000000000000000000000000000300a0ae01000000000000000000000000000000000000000300a2ae01000000000000000000000000000000000000000300a2ae01000000000000000000000000000000000000000300a6ae01000000000000000000000000000000000000000300a6ae01000000000000000000000000000000000000000300aeae01000000000000000000000000000000000000000300aeae01000000000000000000000000000000000000000300b4ae01000000000000000000000000000000000000000300b4ae01000000000000000000000000000000000000000300b8ae01000000000000000000000000000000000000000300c0ae01000000000000000000000000000000000000000300c4ae01000000000000000000000000000000000000000300d0ae01000000000000000000000000000000000000000300d0ae01000000000000000000000000000000000000000300d6ae01000000000000000000000000000000000000000300d6ae01000000000000000000000000000000000000000300daae01000000000000000000000000000000000000000300e2ae01000000000000000000000000000000000000000300e8ae01000000000000000000000000000000000000000300f0ae01000000000000000000000000000000000000000300f4ae0100000000000000000000000000000000000000030000af0100000000000000000000000000000000000000030006af010000000000000000000000000000000000000003000eaf0100000000000000000000000000000000000000030014af010000000000000000000000000000000000000003001caf0100000000000000000000000000000000000000030022af010000000000000000000000000000000000000003002aaf010000000000000000000000000000000000000003002eaf0100000000000000000000000000000000000000030038af0100000000000000000000000000000000000000030038af0100000000000000000000000000000000000000030042af0100000000000000000000000000000000000000030042af0100000000000000000000000000000000000000030044af0100000000000000000000000000000000000000030048af0100000000000000000000000000000000000000030048af0100000000000000000000000000393b00000200030048af0100000000003a00000000000000000000000000030048af0100000000000000000000000000000000000000030048af0100000000000000000000000000000000000000030048af010000000000000000000000000000000000000003004aaf010000000000000000000000000000000000000003004aaf010000000000000000000000000000000000000003004caf01000000000000000000000000008f3b00000000030068af0100000000000000000000000000000000000000030068af0100000000000000000000000000000000000000030068af010000000000000000000000000000000000000003007caf010000000000000000000000000000000000000003007caf010000000000000000000000000000000000000003007eaf0100000000000000000000000000000000000000030082af0100000000000000000000000000000000000000030082af01000000000000000000000000009d3b00000200030082af0100000000002001000000000000000000000000030082af0100000000000000000000000000000000000000030082af0100000000000000000000000000000000000000030082af0100000000000000000000000000000000000000030084af0100000000000000000000000000000000000000030092af0100000000000000000000000000000000000000030094af0100000000000000000000000000000000000000030098af0100000000000000000000000000000000000000030098af010000000000000000000000000000000000000003009aaf010000000000000000000000000000000000000003009aaf01000000000000000000000000000000000000000300a2af01000000000000000000000000000000000000000300a6af01000000000000000000000000000000000000000300a6af01000000000000000000000000000000000000000300aaaf01000000000000000000000000000000000000000300aaaf01000000000000000000000000000000000000000300aeaf01000000000000000000000000000000000000000300aeaf01000000000000000000000000000000000000000300b2af01000000000000000000000000000000000000000300b2af01000000000000000000000000000000000000000300b6af01000000000000000000000000000000000000000300b6af01000000000000000000000000000000000000000300b8af01000000000000000000000000000000000000000300bcaf0100000000000000000000000000d93b000000000300c0af0100000000000000000000000000e73b000001000100ae0501000000000002000000000000000000000000000300c0af01000000000000000000000000000000000000000300caaf01000000000000000000000000000000000000000300ceaf01000000000000000000000000000000000000000300ceaf0100000000000000000000000000133c000000000300d8af0100000000000000000000000000213c000001000100b00501000000000002000000000000000000000000000300e4af01000000000000000000000000000000000000000300e4af01000000000000000000000000000000000000000300e6af01000000000000000000000000004d3c000000000300ecaf01000000000000000000000000005b3c000001000100b20501000000000001000000000000000000000000000300f4af01000000000000000000000000000000000000000300f4af01000000000000000000000000000000000000000300feaf01000000000000000000000000000000000000000300feaf0100000000000000000000000000000000000000030000b00100000000000000000000000000000000000000030000b00100000000000000000000000000000000000000030004b00100000000000000000000000000000000000000030004b00100000000000000000000000000000000000000030006b00100000000000000000000000000000000000000030006b00100000000000000000000000000000000000000030012b00100000000000000000000000000000000000000030012b00100000000000000000000000000000000000000030016b00100000000000000000000000000000000000000030016b00100000000000000000000000000000000000000030018b0010000000000000000000000000000000000000003001cb0010000000000000000000000000000000000000003001cb00100000000000000000000000000000000000000030024b00100000000000000000000000000000000000000030024b0010000000000000000000000000000000000000003002eb0010000000000000000000000000000000000000003002eb00100000000000000000000000000000000000000030032b00100000000000000000000000000000000000000030036b0010000000000000000000000000000000000000003003eb00100000000000000000000000000000000000000030046b0010000000000000000000000000000000000000003005ab0010000000000000000000000000000000000000003005ab0010000000000000000000000000000000000000003005eb00100000000000000000000000000873c0000000003005eb00100000000000000000000000000953c0000010001007005010000000000300000000000000000000000000003005eb00100000000000000000000000000000000000000030068b00100000000000000000000000000000000000000030068b00100000000000000000000000000000000000000030070b00100000000000000000000000000000000000000030070b00100000000000000000000000000c13c00000000030076b00100000000000000000000000000cf3c000001000100ac050100000000000200000000000000000000000000030082b00100000000000000000000000000000000000000030082b00100000000000000000000000000000000000000030084b00100000000000000000000000000000000000000030084b00100000000000000000000000000000000000000030088b0010000000000000000000000000000000000000003008eb0010000000000000000000000000000000000000003009eb001000000000000000000000000000000000000000300a2b001000000000000000000000000000000000000000300a2b00100000000000000000000000000fb3c000002000300a2b001000000000000010000000000000000000000000300a2b001000000000000000000000000000000000000000300a2b001000000000000000000000000000000000000000300a2b001000000000000000000000000000000000000000300a4b001000000000000000000000000000000000000000300b2b001000000000000000000000000000000000000000300b4b001000000000000000000000000000000000000000300b4b001000000000000000000000000000000000000000300bcb001000000000000000000000000000000000000000300bcb001000000000000000000000000000000000000000300beb001000000000000000000000000000000000000000300beb001000000000000000000000000000000000000000300c2b001000000000000000000000000000000000000000300c6b001000000000000000000000000000000000000000300c6b001000000000000000000000000000000000000000300d6b001000000000000000000000000000000000000000300dab001000000000000000000000000000000000000000300deb001000000000000000000000000000000000000000300deb001000000000000000000000000000000000000000300e2b001000000000000000000000000000000000000000300e2b001000000000000000000000000000000000000000300e6b001000000000000000000000000000000000000000300e6b001000000000000000000000000000000000000000300eab001000000000000000000000000000000000000000300eab001000000000000000000000000000000000000000300eeb001000000000000000000000000000000000000000300eeb001000000000000000000000000000000000000000300f0b001000000000000000000000000000000000000000300f2b001000000000000000000000000000000000000000300f2b00100000000000000000000000000343d000000000300fcb0010000000000000000000000000000000000000003000ab1010000000000000000000000000000000000000003000ab1010000000000000000000000000000000000000003000cb10100000000000000000000000000000000000000030016b10100000000000000000000000000000000000000030018b10100000000000000000000000000000000000000030018b10100000000000000000000000000423d00000000030022b10100000000000000000000000000503d000001000100b4050100000000000100000000000000000000000000030030b10100000000000000000000000000000000000000030030b10100000000000000000000000000000000000000030032b10100000000000000000000000000000000000000030032b10100000000000000000000000000000000000000030036b10100000000000000000000000000000000000000030036b10100000000000000000000000000000000000000030038b1010000000000000000000000000000000000000003003cb1010000000000000000000000000000000000000003003cb10100000000000000000000000000000000000000030044b10100000000000000000000000000000000000000030044b1010000000000000000000000000000000000000003004eb1010000000000000000000000000000000000000003004eb10100000000000000000000000000000000000000030052b10100000000000000000000000000000000000000030056b1010000000000000000000000000000000000000003005eb10100000000000000000000000000000000000000030066b101000000000000000000000000007c3d0000000003007ab10100000000000000000000000000000000000000030084b10100000000000000000000000000000000000000030084b1010000000000000000000000000000000000000003008cb1010000000000000000000000000000000000000003008cb101000000000000000000000000008a3d00000000030092b101000000000000000000000000000000000000000300a2b101000000000000000000000000000000000000000300a2b101000000000000000000000000000000000000000300a2b101000000000000000000000000000000000000000300a2b101000000000000000000000000000000000000000300a2b101000000000000000000000000000000000000000300a2b101000000000000000000000000000000000000000300a4b101000000000000000000000000000000000000000300acb101000000000000000000000000000000000000000300aeb101000000000000000000000000000000000000000300aeb101000000000000000000000000000000000000000300bab101000000000000000000000000000000000000000300bab101000000000000000000000000000000000000000300c6b101000000000000000000000000000000000000000300c6b101000000000000000000000000000000000000000300d4b101000000000000000000000000000000000000000300d4b101000000000000000000000000000000000000000300d6b101000000000000000000000000000000000000000300dab101000000000000000000000000000000000000000300dcb101000000000000000000000000000000000000000300deb101000000000000000000000000000000000000000300deb101000000000000000000000000000000000000000300e0b101000000000000000000000000000000000000000300e0b101000000000000000000000000000000000000000300eab101000000000000000000000000000000000000000300ecb101000000000000000000000000000000000000000300f4b101000000000000000000000000000000000000000300f4b101000000000000000000000000000000000000000300fab101000000000000000000000000000000000000000300fab101000000000000000000000000000000000000000300fcb101000000000000000000000000000000000000000300fcb10100000000000000000000000000983d00000000030002b20100000000000000000000000000a63d000001000100b3050100000000000100000000000000000000000000030010b20100000000000000000000000000000000000000030010b20100000000000000000000000000000000000000030012b20100000000000000000000000000000000000000030012b20100000000000000000000000000d23d00000000030018b20100000000000000000000000000e03d00000100010052050100000000000100000000000000000000000000030028b20100000000000000000000000000000000000000030028b2010000000000000000000000000000000000000003002cb2010000000000000000000000000000000000000003002cb20100000000000000000000000000000000000000030036b2010000000000000000000000000000000000000003003ab2010000000000000000000000000000000000000003003ab2010000000000000000000000000000000000000003003ab2010000000000000000000000000000000000000003003ab2010000000000000000000000000000000000000003003ab2010000000000000000000000000000000000000003003cb2010000000000000000000000000000000000000003003cb2010000000000000000000000000000000000000003003eb20100000000000000000000000000000000000000030048b20100000000000000000000000000000000000000030048b201000000000000000000000000000c3e00000200030048b20100000000007200000000000000000000000000030048b20100000000000000000000000000000000000000030048b20100000000000000000000000000000000000000030048b2010000000000000000000000000000000000000003004ab2010000000000000000000000000000000000000003004cb2010000000000000000000000000000000000000003004eb2010000000000000000000000000000000000000003004eb20100000000000000000000000000000000000000030056b20100000000000000000000000000000000000000030056b20100000000000000000000000000000000000000030062b20100000000000000000000000000000000000000030062b20100000000000000000000000000000000000000030064b20100000000000000000000000000000000000000030064b20100000000000000000000000000000000000000030068b20100000000000000000000000000000000000000030068b20100000000000000000000000000000000000000030070b20100000000000000000000000000000000000000030070b20100000000000000000000000000000000000000030078b20100000000000000000000000000000000000000030078b2010000000000000000000000000000000000000003007cb2010000000000000000000000000000000000000003007cb20100000000000000000000000000000000000000030086b20100000000000000000000000000000000000000030086b20100000000000000000000000000000000000000030090b201000000000000000000000000006b3e00000000030090b20100000000000000000000000000000000000000030090b201000000000000000000000000000000000000000300a6b201000000000000000000000000000000000000000300a6b201000000000000000000000000000000000000000300a8b201000000000000000000000000000000000000000300acb201000000000000000000000000000000000000000300acb201000000000000000000000000000000000000000300bab201000000000000000000000000000000000000000300bab201000000000000000000000000000000000000000300bab20100000000000000000000000000793e000002000300bab201000000000072000000000000000000000000000300bab201000000000000000000000000000000000000000300bab201000000000000000000000000000000000000000300bab201000000000000000000000000000000000000000300bcb201000000000000000000000000000000000000000300beb201000000000000000000000000000000000000000300c0b201000000000000000000000000000000000000000300c0b201000000000000000000000000000000000000000300c8b201000000000000000000000000000000000000000300c8b201000000000000000000000000000000000000000300d4b201000000000000000000000000000000000000000300d4b201000000000000000000000000000000000000000300d6b201000000000000000000000000000000000000000300d6b201000000000000000000000000000000000000000300dab201000000000000000000000000000000000000000300dab201000000000000000000000000000000000000000300e2b201000000000000000000000000000000000000000300e2b201000000000000000000000000000000000000000300eab201000000000000000000000000000000000000000300eab201000000000000000000000000000000000000000300eeb201000000000000000000000000000000000000000300eeb201000000000000000000000000000000000000000300f8b201000000000000000000000000000000000000000300f8b20100000000000000000000000000000000000000030002b30100000000000000000000000000d83e00000000030002b30100000000000000000000000000000000000000030002b30100000000000000000000000000000000000000030018b30100000000000000000000000000000000000000030018b3010000000000000000000000000000000000000003001ab3010000000000000000000000000000000000000003001eb3010000000000000000000000000000000000000003001eb3010000000000000000000000000000000000000003002cb3010000000000000000000000000000000000000003002cb3010000000000000000000000000000000000000003002cb30100000000000000000000000000e63e0000020003002cb3010000000000160000000000000000000000000003002cb3010000000000000000000000000000000000000003002cb301000000000000000000000000002e3f0000000003002cb3010000000000000000000000000000000000000003002cb301000000000000000000000000003c3f000001000100b006010000000000020000000000000000000000000003002cb30100000000000000000000000000000000000000030042b30100000000000000000000000000000000000000030042b30100000000000000000000000000000000000000030042b30100000000000000000000000000683f00000200030042b3010000000000a200000000000000000000000000030042b30100000000000000000000000000000000000000030042b30100000000000000000000000000000000000000030042b30100000000000000000000000000000000000000030044b3010000000000000000000000000000000000000003004ab3010000000000000000000000000000000000000003004cb3010000000000000000000000000000000000000003004cb3010000000000000000000000000000000000000003004eb3010000000000000000000000000000000000000003004eb30100000000000000000000000000000000000000030050b30100000000000000000000000000000000000000030050b30100000000000000000000000000c93f00000000030054b30100000000000000000000000000d73f000001000100d8060100000000001100000000000000000000000000030060b30100000000000000000000000000000000000000030060b3010000000000000000000000000000000000000003006cb3010000000000000000000000000003400000000003006cb301000000000000000000000000001140000001000100b806010000000000200000000000000000000000000003006cb30100000000000000000000000000000000000000030080b30100000000000000000000000000000000000000030080b30100000000000000000000000000000000000000030082b30100000000000000000000000000000000000000030086b30100000000000000000000000000000000000000030088b3010000000000000000000000000000000000000003008ab3010000000000000000000000000000000000000003008ab3010000000000000000000000000000000000000003008cb3010000000000000000000000000000000000000003008cb30100000000000000000000000000000000000000030096b30100000000000000000000000000000000000000030098b301000000000000000000000000000000000000000300a0b301000000000000000000000000000000000000000300a0b301000000000000000000000000000000000000000300a6b301000000000000000000000000000000000000000300a6b301000000000000000000000000000000000000000300a8b301000000000000000000000000000000000000000300a8b301000000000000000000000000003d40000000000300aeb301000000000000000000000000000000000000000300bcb301000000000000000000000000000000000000000300bcb301000000000000000000000000000000000000000300beb301000000000000000000000000000000000000000300beb301000000000000000000000000004b40000000000300c4b301000000000000000000000000000000000000000300d4b301000000000000000000000000000000000000000300d4b301000000000000000000000000000000000000000300d8b301000000000000000000000000000000000000000300d8b301000000000000000000000000000000000000000300e0b301000000000000000000000000000000000000000300e4b301000000000000000000000000000000000000000300e4b301000000000000000000000000005940000002000300e4b301000000000070000000000000000000000000000300e4b301000000000000000000000000000000000000000300e4b301000000000000000000000000000000000000000300e4b301000000000000000000000000000000000000000300e6b301000000000000000000000000000000000000000300e8b301000000000000000000000000000000000000000300eab301000000000000000000000000000000000000000300eab301000000000000000000000000000000000000000300f2b301000000000000000000000000000000000000000300f2b301000000000000000000000000000000000000000300fab301000000000000000000000000000000000000000300fab301000000000000000000000000000000000000000300fcb301000000000000000000000000000000000000000300fcb30100000000000000000000000000000000000000030000b40100000000000000000000000000000000000000030000b40100000000000000000000000000000000000000030008b4010000000000000000000000000000000000000003000ab4010000000000000000000000000000000000000003000ab40100000000000000000000000000000000000000030012b40100000000000000000000000000000000000000030012b40100000000000000000000000000000000000000030016b40100000000000000000000000000000000000000030016b40100000000000000000000000000000000000000030020b40100000000000000000000000000000000000000030020b4010000000000000000000000000000000000000003002ab40100000000000000000000000000b9400000000003002ab4010000000000000000000000000000000000000003002ab40100000000000000000000000000000000000000030040b40100000000000000000000000000000000000000030040b40100000000000000000000000000000000000000030042b40100000000000000000000000000000000000000030046b40100000000000000000000000000000000000000030046b40100000000000000000000000000000000000000030054b40100000000000000000000000000000000000000030054b40100000000000000000000000000000000000000030054b40100000000000000000000000000000000000000030054b40100000000000000000000000000000000000000030056b40100000000000000000000000000000000000000030060b40100000000000000000000000000c740000002000300a6b40100000000007c000000000000000000000000000300a6b401000000000000000000000000000000000000000300a6b401000000000000000000000000000000000000000300a8b401000000000000000000000000000000000000000300aeb40100000000000000000000000000000000000000030022b50100000000000000000000000000000000000000030022b50100000000000000000000000000000000000000030024b5010000000000000000000000000000000000000003002cb50100000000000000000000000000000000000000030084b50100000000000000000000000000214100000200030084b50100000000003600000000000000000000000000030084b501000000000000000000000000000000000000000300bab501000000000000000000000000006941000002000300bab501000000000030000000000000000000000000000300bab501000000000000000000000000000000000000000300eab501000000000000000000000000000000000000000300eab501000000000000000000000000000000000000000300ecb501000000000000000000000000000000000000000300f0b50100000000000000000000000000000000000000030036b60100000000000000000000000000b14100000200030036b60100000000008600000000000000000000000000030036b60100000000000000000000000000000000000000030038b60100000000000000000000000000000000000000030044b60100000000000000000000000000104200000000030052b601000000000000000000000000001e420000010001006c0501000000000001000000000000004a420000000003006cb6010000000000000000000000000058420000000003009cb601000000000000000000000000006642000001000100b50501000000000001000000000000000000000000000300bcb601000000000000000000000000009242000002000300bcb601000000000068000000000000000000000000000300bcb601000000000000000000000000000000000000000300beb601000000000000000000000000000000000000000300c8b60100000000000000000000000000d34200000200030024b70100000000007c00000000000000000000000000030024b70100000000000000000000000000000000000000030024b70100000000000000000000000000000000000000030026b7010000000000000000000000000000000000000003002cb701000000000000000000000000002d43000002000300a0b701000000000052000000000000000000000000000300a0b701000000000000000000000000000000000000000300a0b701000000000000000000000000000000000000000300a2b701000000000000000000000000000000000000000300a8b701000000000000000000000000000000000000000300f2b701000000000000000000000000000000000000000300f2b701000000000000000000000000000000000000000300f4b701000000000000000000000000000000000000000300f8b70100000000000000000000000000000000000000030048b80100000000000000000000000000604300000200030048b80100000000008201000000000000000000000000030048b8010000000000000000000000000000000000000003004ab80100000000000000000000000000000000000000030058b8010000000000000000000000000091430000000003002ab901000000000000000000000000009f4300000100010090070100000000001c00000000000000a94300000000030034b90100000000000000000000000000b7430000000003003eb90100000000000000000000000000c54300000000030052b90100000000000000000000000000d3430000000003005ab90100000000000000000000000000e143000001000100100701000000000020000000000000000b4400000000030068b901000000000000000000000000001944000001000100f6070100000000002f00000000000000444400000000030076b901000000000000000000000000005244000001000100250801000000000032000000000000007d4400000000030090b901000000000000000000000000008b4400000000030098b90100000000000000000000000000994400000100010068070100000000002000000000000000c344000000000300b2b90100000000000000000000000000d144000001000100ac070100000000001c00000000000000fc44000000000300bcb901000000000000000000000000000a45000001000100c8070100000000002e000000000000000000000000000300cab901000000000000000000000000003545000002000300cab901000000000028000000000000000000000000000300cab901000000000000000000000000009045000000000300d0b901000000000000000000000000009e45000001000100600d01000000000050000000000000000846000000000300dab901000000000000000000000000001646000001000100b00d01000000000050000000000000000000000000000300f2b901000000000000000000000000000000000000000300f2b901000000000000000000000000000000000000000300f4b90100000000000000000000000000844600000000030014ba0100000000000000000000000000924600000000030020ba0100000000000000000000000000a04600000100010030070100000000001800000000000000ca4600000000030028ba0100000000000000000000000000d8460000010001004807010000000000200000000000000002470000000003003eba0100000000000000000000000000104700000100010057080100000000002600000000000000000000000000030054ba01000000000000000000000000003b4700000200030054ba0100000000006800000000000000000000000000030054ba0100000000000000000000000000000000000000030056ba010000000000000000000000000000000000000003005aba01000000000000000000000000007a4700000000030086ba010000000000000000000000000088470000000003008eba01000000000000000000000000009647000000000300a8ba0100000000000000000000000000a4470000010001007d080100000000000d000000000000000000000000000300bcba01000000000000000000000000000000000000000300bcba01000000000000000000000000000000000000000300beba01000000000000000000000000000000000000000300c0ba0100000000000000000000000000cf47000000000300d8ba0100000000000000000000000000dd470000010001008a080100000000000e000000000000000000000000000300ecba01000000000000000000000000000000000000000300ecba01000000000000000000000000000000000000000300eeba0100000000000000000000000000000000000000030000bb010000000000000000000000000008480000000003007cbb010000000000000000000000000016480000000003000abc0100000000000000000000000000244800000000030014bc010000000000000000000000000032480000000003001ebc0100000000000000000000000000404800000000030028bc01000000000000000000000000004e4800000000030032bc01000000000000000000000000005c480000000003003cbc0100000000000000000000000000000000000000030052bc0100000000000000000000000000000000000000030052bc0100000000000000000000000000000000000000030054bc0100000000000000000000000000000000000000030058bc01000000000000000000000000006a48000000000300a0bc01000000000000000000000000000000000000000300b6bc01000000000000000000000000000000000000000300b6bc01000000000000000000000000000000000000000300b8bc01000000000000000000000000000000000000000300bebc01000000000000000000000000007848000000000300f8bc0100000000000000000000000000864800000000030000bd010000000000000000000000000094480000000003001abd0100000000000000000000000000a24800000100010098080100000000000e0000000000000000000000000003002ebd010000000000000000000000000000000000000003002ebd0100000000000000000000000000000000000000030030bd0100000000000000000000000000000000000000030036bd0100000000000000000000000000cd4800000000030076bd0100000000000000000000000000db480000000003007ebd0100000000000000000000000000e94800000000030098bd0100000000000000000000000000f748000001000100b4080100000000000d000000000000000000000000000300acbd01000000000000000000000000000000000000000300acbd01000000000000000000000000000000000000000300aebd01000000000000000000000000000000000000000300b6bd0100000000000000000000000000224900000000030018be0100000000000000000000000000304900000000030020be01000000000000000000000000003e490000000003003abe01000000000000000000000000004c49000001000100c108010000000000120000000000000000000000000003004ebe010000000000000000000000000077490000020003004ebe0100000000007a0000000000000000000000000003004ebe0100000000000000000000000000000000000000030050be0100000000000000000000000000000000000000030056be0100000000000000000000000000db49000000000300a6be01000000000000000000000000000000000000000300c8be01000000000000000000000000000000000000000300c8be01000000000000000000000000000000000000000300cabe01000000000000000000000000000000000000000300d6be0100000000000000000000000000e94900000000030030bf0100000000000000000000000000f749000001000100d808010000000000200000000000000000000000000003007abf0100000000000000000000000000224a0000020003007abf010000000000100000000000000000000000000003007abf010000000000000000000000000000000000000003008abf0100000000000000000000000000734a0000020003008abf0100000000008c0000000000000000000000000003008abf010000000000000000000000000000000000000003008cbf0100000000000000000000000000000000000000030094bf0100000000000000000000000000000000000000030016c00100000000000000000000000000b64a00000200030016c00100000000004a00000000000000000000000000030016c00100000000000000000000000000000000000000030060c001000000000000000000000000001a4b00000200030060c00100000000007200000000000000000000000000030060c00100000000000000000000000000000000000000030062c0010000000000000000000000000000000000000003006ac001000000000000000000000000009b4b000000000300b4c00100000000000000000000000000a94b000001000100a0090100000000001c000000000000000000000000000300d2c001000000000000000000000000000000000000000300d2c00100000000000000000000000000b34b00000000030072c10100000000000000000000000000c14b00000000030088c10100000000000000000000000000000000000000030092c10100000000000000000000000000cf4b00000200030092c10100000000002400000000000000000000000000030092c10100000000000000000000000000000000000000030094c10100000000000000000000000000000000000000030096c101000000000000000000000000000000000000000300b6c10100000000000000000000000000144c000002000300b6c101000000000024000000000000000000000000000300b6c101000000000000000000000000000000000000000300b8c101000000000000000000000000000000000000000300bac101000000000000000000000000000000000000000300dac10100000000000000000000000000594c000002000300dac101000000000014010000000000000000000000000300dac101000000000000000000000000000000000000000300dcc101000000000000000000000000000000000000000300f4c101000000000000000000000000000000000000000300eec20100000000000000000000000000744d000002000300eec20100000000006c000000000000000000000000000300eec2010000000000000000000000000000000000000003005ac30100000000000000000000000000194e0000020003005ac30100000000007e0300000000000000000000000003005ac3010000000000000000000000000000000000000003005cc30100000000000000000000000000000000000000030076c30100000000000000000000000000674f00000200030046ca010000000000e802000000000000d74f00000200030040c701000000000006030000000000003e500000020003002ecd010000000000d002000000000000a450000002000300fecf010000000000ae020000000000000000000000000300d8c601000000000000000000000000000000000000000300d8c60100000000000000000000000000000000000000030040c70100000000000000000000000000000000000000030040c70100000000000000000000000000000000000000030042c7010000000000000000000000000000000000000003005cc70100000000000000000000000000025100000000030002ca010000000000000000000000000010510000010001002e0b0100000000001b000000000000003b510000000003000eca010000000000000000000000000049510000000003001cca0100000000000000000000000000575100000000030026ca0100000000000000000000000000655100000000030030ca0100000000000000000000000000000000000000030046ca0100000000000000000000000000000000000000030046ca0100000000000000000000000000000000000000030048ca0100000000000000000000000000000000000000030062ca010000000000000000000000000073510000000003000acd0100000000000000000000000000815100000000030018cd010000000000000000000000000000000000000003002ecd010000000000000000000000000000000000000003002ecd0100000000000000000000000000000000000000030030cd010000000000000000000000000000000000000003004acd01000000000000000000000000008f51000000000300b6cf01000000000000000000000000009d51000000000300c2cf0100000000000000000000000000ab51000000000300d0cf0100000000000000000000000000b951000000000300decf0100000000000000000000000000c751000000000300e8cf01000000000000000000000000000000000000000300fecf01000000000000000000000000000000000000000300fecf0100000000000000000000000000000000000000030000d0010000000000000000000000000000000000000003001ad00100000000000000000000000000d55100000000030096d201000000000000000000000000000000000000000300acd20100000000000000000000000000e351000002000300acd201000000000024000000000000000000000000000300acd201000000000000000000000000000000000000000300aed201000000000000000000000000000000000000000300b0d201000000000000000000000000000000000000000300d0d201000000000000000000000000002852000002000300d0d201000000000024000000000000000000000000000300d0d201000000000000000000000000000000000000000300d2d201000000000000000000000000000000000000000300d4d201000000000000000000000000000000000000000300f4d201000000000000000000000000006d52000002000300f4d201000000000028010000000000000000000000000300f4d201000000000000000000000000000000000000000300f6d2010000000000000000000000000000000000000003000cd3010000000000000000000000000000000000000003001cd4010000000000000000000000000088530000020003001cd4010000000000680000000000000000000000000003001cd4010000000000000000000000000000000000000003001ed4010000000000000000000000000000000000000003002cd40100000000000000000000000000000000000000030084d401000000000000000000000000002d5400000200030084d40100000000000403000000000000000000000000030084d40100000000000000000000000000000000000000030088d401000000000000000000000000000000000000000300bcd401000000000000000000000000007b5500000200030088d701000000000066000000000000004356000002000300b4da0100000000004602000000000000b356000002000300eed7010000000000c6020000000000001a57000002000300fadc0100000000008e02000000000000805700000200030088df0100000000000202000000000000000000000000030088d70100000000000000000000000000000000000000030088d701000000000000000000000000000000000000000300eed701000000000000000000000000000000000000000300eed701000000000000000000000000000000000000000300f2d70100000000000000000000000000000000000000030026d80100000000000000000000000000de5700000000030070da0100000000000000000000000000ec570000000003007cda0100000000000000000000000000fa570000000003008ada0100000000000000000000000000085800000000030094da010000000000000000000000000016580000000003009eda01000000000000000000000000000000000000000300b4da01000000000000000000000000000000000000000300b4da01000000000000000000000000000000000000000300b6da01000000000000000000000000000000000000000300d0da01000000000000000000000000002458000000000300d6dc01000000000000000000000000003258000000000300e4dc01000000000000000000000000000000000000000300fadc01000000000000000000000000000000000000000300fadc01000000000000000000000000000000000000000300fedc0100000000000000000000000000000000000000030032dd0100000000000000000000000000405800000000030040df01000000000000000000000000004e580000000003004cdf01000000000000000000000000005c580000000003005adf01000000000000000000000000006a5800000000030068df0100000000000000000000000000785800000000030072df0100000000000000000000000000000000000000030088df0100000000000000000000000000000000000000030088df010000000000000000000000000000000000000003008adf01000000000000000000000000000000000000000300a4df0100000000000000000000000000865800000000030074e1010000000000000000000000000000000000000003008ae1010000000000000000000000000094580000020003008ae1010000000000362900000000000000000000000003008ae1010000000000000000000000000000000000000003008ee101000000000000000000000000000000000000000300b8e10100000000000000000000000000c458000002000300621002000000000006040000000000000759000002000300501e02000000000050010000000000003f59000002000300a01f0200000000000c030000000000007f590000020003006814020000000000e8090000000000000000000000000300c00a0200000000000000000000000000b059000000000400a09a0200000000000000000000000000bb59000002000300c00a0200000000008c000000000000000000000000000300c00a02000000000000000000000000000000000000000300c20a02000000000000000000000000000000000000000300c80a0200000000000000000000000000085a000000000300e20a020000000000000000000000000000000000000003004c0b0200000000000000000000000000165a0000020003004c0b020000000000cc0100000000000000000000000003004c0b02000000000000000000000000000000000000000300500b02000000000000000000000000000000000000000300680b02000000000000000000000000004e5a000000000300820b02000000000000000000000000005c5a00000200030074260200000000006a000000000000008a5a000002000300180d020000000000f600000000000000cd5a000000000300720c0200000000000000000000000000db5a000000000300960c0200000000000000000000000000e95a0000020003000e0e02000000000054020000000000000000000000000300180d02000000000000000000000000000000000000000300180d020000000000000000000000000000000000000003001c0d02000000000000000000000000000000000000000300300d020000000000000000000000000000000000000003000e0e020000000000000000000000000000000000000003000e0e02000000000000000000000000000000000000000300120e020000000000000000000000000000000000000003002a0e020000000000000000000000000000000000000003006210020000000000000000000000000000000000000003006210020000000000000000000000000000000000000003006410020000000000000000000000000000000000000003007a1002000000000000000000000000002c5b000000000300521402000000000000000000000000003a5b000001000100c0090100000000002e0000000000000000000000000003006814020000000000000000000000000000000000000003006814020000000000000000000000000000000000000003006a1402000000000000000000000000000000000000000300821402000000000000000000000000000000000000000300501e0200000000000000000000000000655b000000000400a89a0200000000000000000000000000705b000000000400b09a02000000000000000000000000007b5b000000000400b89a0200000000000000000000000000865b000000000400c09a02000000000000000000000000000000000000000300501e02000000000000000000000000000000000000000300521e02000000000000000000000000000000000000000300641e0200000000000000000000000000915b000000000300901e02000000000000000000000000009f5b000000000300981e0200000000000000000000000000ad5b000000000300b21e0200000000000000000000000000bb5b000000000300ba1e0200000000000000000000000000c95b0000000003008c1f02000000000000000000000000000000000000000300a01f02000000000000000000000000000000000000000300a01f02000000000000000000000000000000000000000300a21f02000000000000000000000000000000000000000300bc1f0200000000000000000000000000d75b000002000300ac22020000000000c8030000000000000000000000000300ac2202000000000000000000000000000000000000000300ac2202000000000000000000000000000000000000000300ae2202000000000000000000000000000000000000000300be22020000000000000000000000000000000000000003007426020000000000000000000000000000000000000003007426020000000000000000000000000000000000000003007626020000000000000000000000000000000000000003007e2602000000000000000000000000001b5c000000000300a62602000000000000000000000000000000000000000300de260200000000000000000000000000295c000000000400c89a0200000000000000000000000000345c000002000300de260200000000008c000000000000000000000000000300de2602000000000000000000000000000000000000000300e02602000000000000000000000000000000000000000300e6260200000000000000000000000000815c0000000003000027020000000000000000000000000000000000000003006a2702000000000000000000000000008f5c0000020003006a27020000000000720000000000000000000000000003006a27020000000000000000000000000000000000000003006c270200000000000000000000000000000000000000030074270200000000000000000000000000105d000000000300c82702000000000000000000000000000000000000000300dc2702000000000000000000000000000000000000000300dc2702000000000000000000000000000000000000000300e02702000000000000000000000000000000000000000300f82702000000000000000000000000001e5d000002000300aa2a0200000000003200000000000000905d000000000300f22902000000000000000000000000009e5d0000000003008a2a0200000000000000000000000000ac5d000000000300922a0200000000000000000000000000ba5d000001000100600a01000000000020000000000000000000000000000300aa2a02000000000000000000000000000000000000000300aa2a02000000000000000000000000000000000000000300ac2a02000000000000000000000000000000000000000300b02a02000000000000000000000000000000000000000300dc2a02000000000000000000000000000000000000000300dc2a02000000000000000000000000000000000000000300de2a02000000000000000000000000000000000000000300f42a0200000000000000000000000000e55d000000000300b22d0200000000000000000000000000f35d000000000300c62d0200000000000000000000000000015e000001000100e00c0100000000002b000000000000002d5e000000000300d42d02000000000000000000000000003b5e000000000300dc2d02000000000000000000000000000000000000000300f42d02000000000000000000000000000000000000000300f42d02000000000000000000000000000000000000000300f62d02000000000000000000000000000000000000000300102e0200000000000000000000000000495e0000000003003e310200000000000000000000000000575e00000000030052310200000000000000000000000000655e0000000003005a310200000000000000000000000000735e000001000100200a01000000000020000000000000009e5e00000000030072310200000000000000000000000000ac5e0000010001000b0d010000000000290000000000000000000000000003008031020000000000000000000000000000000000000003008031020000000000000000000000000000000000000003008231020000000000000000000000000000000000000003009c310200000000000000000000000000d85e000000000300ce340200000000000000000000000000e65e000000000300e2340200000000000000000000000000f45e000000000300ea340200000000000000000000000000025f00000000030002350200000000000000000000000000105f000001000100340d0100000000002c0000000000000000000000000003001035020000000000000000000000000000000000000003001035020000000000000000000000000000000000000003001235020000000000000000000000000000000000000003002c3502000000000000000000000000003c5f000000000300dc3802000000000000000000000000004a5f000000000300f0380200000000000000000000000000585f000000000300f8380200000000000000000000000000665f00000000030008390200000000000000000000000000745f00000000030010390200000000000000000000000000825f00000000030020390200000000000000000000000000905f000000000300283902000000000000000000000000009e5f00000000030032390200000000000000000000000000ac5f0000000003003a39020000000000000000000000000000000000000003005e39020000000000000000000000000000000000000003005e39020000000000000000000000000000000000000003006039020000000000000000000000000000000000000003006c390200000000000000000000000000ba5f000000000300be3a02000000000000000000000000000000000000000300e43a02000000000000000000000000000000000000000300e43a02000000000000000000000000000000000000000300e63a02000000000000000000000000000000000000000300003b0200000000000000000000000000c85f000000000300063d0200000000000000000000000000d65f0000000003001a3d0200000000000000000000000000e45f000000000300223d020000000000000000000000000000000000000003003a3d020000000000000000000000000000000000000003003a3d020000000000000000000000000000000000000003003c3d02000000000000000000000000000000000000000300423d0200000000000000000000000000f25f0000000003003a3e02000000000000000000000000000060000000000300423e02000000000000000000000000000e600000000003004c3e02000000000000000000000000001c60000000000300543e02000000000000000000000000002a60000000000300643e020000000000000000000000000038600000000003006c3e020000000000000000000000000046600000000003007c3e02000000000000000000000000005460000000000300843e020000000000000000000000000062600000000003009e3e02000000000000000000000000007060000001000100a6080100000000000e000000000000000000000000000300b23e02000000000000000000000000000000000000000300b23e02000000000000000000000000000000000000000300b43e02000000000000000000000000000000000000000300ce3e02000000000000000000000000009b60000000000300c4400200000000000000000000000000a960000000000300d8400200000000000000000000000000b760000000000300e0400200000000000000000000000000c560000000000300f840020000000000000000000000000000000000000003000641020000000000000000000000000000000000000003000641020000000000000000000000000000000000000003000a41020000000000000000000000000000000000000003003e410200000000000000000000000000d3600000000003006c470200000000000000000000000000e1600000000003002e480200000000000000000000000000ef6000000100010080020100000000001c00000000000000f5600000000003004c4802000000000000000000000000000361000000000300544802000000000000000000000000001161000001000100400a010000000000200000000000000000000000000003006c48020000000000000000000000000000000000000003006c48020000000000000000000000000000000000000003007048020000000000000000000000000000000000000003007c4802000000000000000000000000000000000000000300e04802000000000000000000000000000000000000000300e04802000000000000000000000000000000000000000300e448020000000000000000000000000000000000000003001849020000000000000000000000000000000000000003001849020000000000000000000000000000000000000003001a4902000000000000000000000000003c61000000000300744a02000000000000000000000000004a610000000003002e6402000000000000000000000000005861000000000300506402000000000000000000000000006661000000000300ba7602000000000000000000000000007461000000000100b00101000000000000000000000000007f61000000000300988102000000000000000000000000008b61000000000300ee7602000000000000000000000000009761000000000300c2780200000000000000000000000000a361000000000300267b0200000000000000000000000000af61000000000300e27c0200000000000000000000000000bb61000000000300327d0200000000000000000000000000c761000000000300b0810200000000000000000000000000d561000000000300c2810200000000000000000000000000e361000000000300d0810200000000000000000000000000f161000000000300de810200000000000000000000000000ff61000000000300e88102000000000000000000000000000d62000000000300f28102000000000000000000000000001b62000000000300fc81020000000000000000000000000029620000000003001682020000000000000000000000000037620000000003002c8202000000000000000000000000004562000000000300368202000000000000000000000000005362000000000300448202000000000000000000000000006162000000000300588202000000000000000000000000006f62000000000300628202000000000000000000000000007d620000000003006c8202000000000000000000000000008b6200000000030076820200000000000000000000000000996200000000030080820200000000000000000000000000a7620000000003008a820200000000000000000000000000b5620000000003009e820200000000000000000000000000c362000000000300a8820200000000000000000000000000d162000000000300b2820200000000000000000000000000df62000000000300bc820200000000000000000000000000ed62000000000300c6820200000000000000000000000000fb62000000000300d08202000000000000000000000000000963000000000300ee8202000000000000000000000000001763000000000300f882020000000000000000000000000025630000000003000283020000000000000000000000000033630000000003001283020000000000000000000000000041630000000003001c8302000000000000000000000000000000000000000300268302000000000000000000000000004f63000001000600889b02000000000000100800000000007e6300000100060088ab0a00000000000010000000000000b363000001000100dc030100000000002300000000000000de63000001000100100401000000000033000000000000000964000001000100f8080100000000000a00000000000000346400000100010002090100000000000a000000000000005f640000010001000c090100000000000b000000000000008a6400000100010017090100000000000600000000000000b5640000010001001d090100000000000600000000000000e064000001000100230901000000000009000000000000000b650000010001002c0901000000000006000000000000000000000000000800000000000000000000000000000000000000000000000b009c2b00000000000000000000000000000000000000000b00234600000000000000000000000000003665000000000f00000000000000000000000000000000000000000000000b00521300000000000000000000000000000000000000000b009b2f00000000000000000000000000000000000000000b00000000000000000000000000000000000000000000000b00494f00000000000000000000000000000000000000000b00503800000000000000000000000000000000000000000800510000000000000000000000000000000000000000000b00811700000000000000000000000000004a65000000000f005c0000000000000000000000000000000000000000000a00701100000000000000000000000000000000000000000b00621a00000000000000000000000000000000000000000b00840500000000000000000000000000000000000000000b002f0d00000000000000000000000000000000000000000b00b71700000000000000000000000000000000000000000b00c83500000000000000000000000000000000000000000b00dd0c00000000000000000000000000000000000000000b00813f00000000000000000000000000000000000000000b00833300000000000000000000000000000000000000000b00d23800000000000000000000000000000000000000000b003f2500000000000000000000000000000000000000000b00cb2a00000000000000000000000000000000000000000b00932300000000000000000000000000000000000000000b00122d00000000000000000000000000000000000000000b00944900000000000000000000000000000000000000000b00a63b00000000000000000000000000000000000000000b005b3a00000000000000000000000000000000000000000b00770c00000000000000000000000000000000000000000b00f90300000000000000000000000000000000000000000b005f0d00000000000000000000000000000000000000000b00844200000000000000000000000000000000000000000b009c3300000000000000000000000000000000000000000b00b41800000000000000000000000000000000000000000b00ff0b00000000000000000000000000000000000000000b00c13700000000000000000000000000000000000000000b00a60000000000000000000000000000000000000000000b003c4a00000000000000000000000000000000000000000b00241400000000000000000000000000000000000000000b002d4400000000000000000000000000000000000000000b00e74800000000000000000000000000000000000000000b00900500000000000000000000000000000000000000000b00b80800000000000000000000000000000000000000000b00cc0000000000000000000000000000000000000000000b003c2a00000000000000000000000000000000000000000b007f3300000000000000000000000000000000000000000b00821300000000000000000000000000000000000000000b007c3400000000000000000000000000000000000000000b00ca4b00000000000000000000000000000000000000000b007b2900000000000000000000000000000000000000000b00514100000000000000000000000000000000000000000b005d1400000000000000000000000000000000000000000b008b4900000000000000000000000000000000000000000b007b3e00000000000000000000000000000000000000000b00214c00000000000000000000000000000000000000000b00763100000000000000000000000000000000000000000b00231700000000000000000000000000000000000000000b00623800000000000000000000000000000000000000000a00000000000000000000000000000000000000000000000a00400000000000000000000000000000000000000000000a00700000000000000000000000000000000000000000000a00a00000000000000000000000000000000000000000000b00550c00000000000000000000000000000000000000000b006e2d00000000000000000000000000000000000000000b00ac3e00000000000000000000000000000000000000000b006b1b00000000000000000000000000000000000000000b00f20400000000000000000000000000000000000000000b00e81600000000000000000000000000000000000000000b00db1000000000000000000000000000000000000000000b00d13000000000000000000000000000000000000000000b00752b00000000000000000000000000000000000000000b00512b00000000000000000000000000000000000000000b00281500000000000000000000000000000000000000000b007f1d00000000000000000000000000000000000000000b004e4700000000000000000000000000000000000000000b00884a00000000000000000000000000000000000000000b00093c00000000000000000000000000000000000000000b009d1500000000000000000000000000000000000000000b00163100000000000000000000000000000000000000000a00200900000000000000000000000000000000000000000a00500900000000000000000000000000000000000000000a00800900000000000000000000000000000000000000000a00b00900000000000000000000000000000000000000000a00e00900000000000000000000000000000000000000000b00c60700000000000000000000000000000000000000000b005f3500000000000000000000000000000000000000000b000f0f00000000000000000000000000000000000000000b001c2900000000000000000000000000000000000000000a00100e00000000000000000000000000000000000000000a00400e00000000000000000000000000000000000000000a00700e00000000000000000000000000000000000000000a00a00e00000000000000000000000000000000000000000a00d00e00000000000000000000000000000000000000000b000e4800000000000000000000000000000000000000000b00724800000000000000000000000000000000000000000a00000f00000000000000000000000000000000000000000a00300f00000000000000000000000000000000000000000a00600f00000000000000000000000000000000000000000a00900f00000000000000000000000000000000000000000a00c00f00000000000000000000000000000000000000000b00210800000000000000000000000000000000000000000b001f0300000000000000000000000000000000000000000a00801000000000000000000000000000000000000000000a00b01000000000000000000000000000000000000000000a00e01000000000000000000000000000000000000000000a00101100000000000000000000000000000000000000000a00401100000000000000000000000000000000000000000b00a44d00000000000000000000000000000000000000000b00e90a00000000000000000000000000000000000000000b001e0b00000000000000000000000000000000000000000b007f0300000000000000000000000000000000000000000b007a3100000000000000000000000000000000000000000b00964c00000000000000000000000000000000000000000b00194400000000000000000000000000000000000000000b006b0d00000000000000000000000000000000000000000b00880500000000000000000000000000000000000000000b00890200000000000000000000000000000000000000000b00b83400000000000000000000000000000000000000000a00d00000000000000000000000000000000000000000000a00100100000000000000000000000000000000000000000a00400100000000000000000000000000000000000000000a00700100000000000000000000000000000000000000000a00a00100000000000000000000000000000000000000000a00d00100000000000000000000000000000000000000000a00000200000000000000000000000000000000000000000a00300200000000000000000000000000000000000000000a00800200000000000000000000000000000000000000000b00454b00000000000000000000000000000000000000000b000c3100000000000000000000000000000000000000000a00b00200000000000000000000000000000000000000000a00e00200000000000000000000000000000000000000000a00100300000000000000000000000000000000000000000a00400300000000000000000000000000000000000000000a00700300000000000000000000000000000000000000000a00a00300000000000000000000000000000000000000000a00d00300000000000000000000000000000000000000000a00000400000000000000000000000000000000000000000a00300400000000000000000000000000000000000000000a00800400000000000000000000000000000000000000000a00b00400000000000000000000000000000000000000000a00000500000000000000000000000000000000000000000a00300500000000000000000000000000000000000000000a00800500000000000000000000000000000000000000000a00b00500000000000000000000000000000000000000000a00f00500000000000000000000000000000000000000000a00600600000000000000000000000000000000000000000a00b00600000000000000000000000000000000000000000a00f00600000000000000000000000000000000000000000a00200700000000000000000000000000000000000000000a00500700000000000000000000000000000000000000000b00773b00000000000000000000000000000000000000000b002b3000000000000000000000000000000000000000000b00bf1800000000000000000000000000000000000000000b00642d00000000000000000000000000000000000000000b00fe3300000000000000000000000000000000000000000b00442b00000000000000000000000000000000000000000b00e82800000000000000000000000000000000000000000b00111e00000000000000000000000000000000000000000b00db0700000000000000000000000000000000000000000b00252500000000000000000000000000000000000000000b00ec1b00000000000000000000000000000000000000000b00801800000000000000000000000000000000000000000b000e3200000000000000000000000000000000000000000b00143200000000000000000000000000000000000000000b00544d00000000000000000000000000000000000000000b00a61b00000000000000000000000000000000000000000b00ac0900000000000000000000000000000000000000000b00104d00000000000000000000000000000000000000000b003e1000000000000000000000000000000000000000000b00d10900000000000000000000000000000000000000000b00803c00000000000000000000000000000000000000000a00800700000000000000000000000000000000000000000a00b00700000000000000000000000000000000000000000a00e00700000000000000000000000000000000000000000a00100800000000000000000000000000000000000000000a00400800000000000000000000000000000000000000000a00700800000000000000000000000000000000000000000a00a00800000000000000000000000000000000000000000a00e00800000000000000000000000000000000000000000b00f10100000000000000000000000000000000000000000b00fa3f00000000000000000000000000000000000000000b00f83b00000000000000000000000000000000000000000b00273b00000000000000000000000000000000000000000b006a3800000000000000000000000000000000000000000a00100a00000000000000000000000000000000000000000a00400a00000000000000000000000000000000000000000a00700a00000000000000000000000000000000000000000a00a00a00000000000000000000000000000000000000000a00d00a00000000000000000000000000000000000000000a00000b00000000000000000000000000000000000000000b00874000000000000000000000000000000000000000000b00084800000000000000000000000000000000000000000b00920400000000000000000000000000000000000000000b00641b00000000000000000000000000000000000000000b00ca2400000000000000000000000000000000000000000b006a2b00000000000000000000000000000000000000000b00144d00000000000000000000000000000000000000000b00294a00000000000000000000000000000000000000000b006f0a00000000000000000000000000000000000000000a00b00b00000000000000000000000000000000000000000a00e00b00000000000000000000000000000000000000000a00100c00000000000000000000000000000000000000000a00400c00000000000000000000000000000000000000000a00700c00000000000000000000000000000000000000000a00b00c00000000000000000000000000000000000000000b008b1e00000000000000000000000000000000000000000b00304b00000000000000000000000000000000000000000b00501e00000000000000000000000000000000000000000b00363000000000000000000000000000000000000000000b00a30900000000000000000000000000000000000000000b00f73700000000000000000000000000000000000000000b00591b00000000000000000000000000000000000000000b003b3000000000000000000000000000000000000000000b00ec0400000000000000000000000000000000000000000b00cf0e00000000000000000000000000000000000000000b00de4c00000000000000000000000000000000000000000b00773000000000000000000000000000000000000000000b00c83a00000000000000000000000000000000000000000b004b0500000000000000000000000000000000000000000a00f00c00000000000000000000000000000000000000000a00200d00000000000000000000000000000000000000000a00500d00000000000000000000000000000000000000000a00800d00000000000000000000000000000000000000000a00b00d00000000000000000000000000000000000000000a00e00d00000000000000000000000000000000000000000b00413400000000000000000000000000000000000000000b00ba2400000000000000000000000000000000000000000b00fb3200000000000000000000000000000000000000000a00300b00000000000000000000000000000000000000000b00d51900000000000000000000000000000000000000000b00013300000000000000000000000000000000000000000b00d74700000000000000000000000000000000000000000b001e4f00000000000000000000000000000000000000000b00744b00000000000000000000000000000000000000000b003a4500000000000000000000000000000000000000000b00654500000000000000000000000000000000000000000a00700b00000000000000000000000000000000000000000b00d13a00000000000000000000000000000000000000000b002a0a00000000000000000000000000000000000000000b00011100000000000000000000000000000000000000000b00d30c00000000000000000000000000000000000000000b00373300000000000000000000000000000000000000000b004c1100000000000000000000000000000000000000000b00c73c00000000000000000000000000000000000000000b009b4d00000000000000000000000000000000000000000b001a4c00000000000000000000000000000000000000000b00340a00000000000000000000000000000000000000000b00824f00000000000000000000000000000000000000000b004b2f00000000000000000000000000000000000000000b00d00700000000000000000000000000000000000000000b00512f00000000000000000000000000000000000000000b00d71000000000000000000000000000000000000000000b00872900000000000000000000000000000000000000000b00190f00000000000000000000000000000000000000000b003b4b00000000000000000000000000000000000000000b00541700000000000000000000000000000000000000000b00103100000000000000000000000000000000000000000b00364000000000000000000000000000000000000000000b00301300000000000000000000000000000000000000000b00681000000000000000000000000000000000000000000b00373400000000000000000000000000000000000000000b00cb3c00000000000000000000000000000000000000000b00ab0a00000000000000000000000000000000000000000b00b51100000000000000000000000000000000000000000b00893400000000000000000000000000000000000000000b00c81e00000000000000000000000000000000000000000b00472500000000000000000000000000000000000000000b00523600000000000000000000000000000000000000000b00d14800000000000000000000000000000000000000000b00013e00000000000000000000000000000000000000000b00c10100000000000000000000000000000000000000000b00982c00000000000000000000000000000000000000000b004c4400000000000000000000000000000000000000000b00384e00000000000000000000000000000000000000000b00304100000000000000000000000000000000000000000b00c71c00000000000000000000000000000000000000000b00dc3f00000000000000000000000000000000000000000b00243900000000000000000000000000000000000000000b00120000000000000000000000000000000000000000000b00cb1b00000000000000000000000000000000000000000b00a82f00000000000000000000000000000000000000000b00d64c00000000000000000000000000000000000000000b00cd3400000000000000000000000000000000000000000b00a32300000000000000000000000000000000000000000b00b32300000000000000000000000000000000000000000b00373700000000000000000000000000000000000000000b002e4e00000000000000000000000000000000000000000b00db3900000000000000000000000000000000000000000b00740b00000000000000000000000000000000000000000b00eb3d00000000000000000000000000000000000000000b004d0c00000000000000000000000000000000000000000b00411d00000000000000000000000000000000000000000b00024500000000000000000000000000000000000000000b00b11200000000000000000000000000000000000000000b00f81b00000000000000000000000000000000000000000b00771c00000000000000000000000000000000000000000b002d2a00000000000000000000000000000000000000000b00034700000000000000000000000000000000000000000b005d4a00000000000000000000000000000000000000000b00532700000000000000000000000000000000000000000b00d14000000000000000000000000000000000000000000b00180600000000000000000000000000000000000000000b00e84000000000000000000000000000000000000000000b00684400000000000000000000000000000000000000000b00620900000000000000000000000000000000000000000b006b2a00000000000000000000000000000000000000000b00b72a00000000000000000000000000000000000000000b00303b00000000000000000000000000000000000000000b00da3d00000000000000000000000000000000000000000b00db1a00000000000000000000000000000000000000000b00f81200000000000000000000000000000000000000000b00bc4400000000000000000000000000000000000000000b00563200000000000000000000000000000000000000000b00ed2700000000000000000000000000000000000000000b00da0900000000000000000000000000000000000000000b005b0e00000000000000000000000000000000000000000b00521900000000000000000000000000000000000000000b004c0400000000000000000000000000000000000000000b00311b00000000000000000000000000000000000000000b00b60700000000000000000000000000000000000000000b00bd4500000000000000000000000000000000000000000b00b53c00000000000000000000000000000000000000000b00b40300000000000000000000000000000000000000000b00af0500000000000000000000000000000000000000000b00c53400000000000000000000000000000000000000000b004d3700000000000000000000000000000000000000000b001d2b00000000000000000000000000000000000000000b00f20d00000000000000000000000000000000000000000b00261300000000000000000000000000000000000000000b005a4100000000000000000000000000000000000000000b00ea3300000000000000000000000000000000000000000b00653a00000000000000000000000000000000000000000b00fa0100000000000000000000000000000000000000000b00b14900000000000000000000000000000000000000000b00673200000000000000000000000000000000000000000b00f41800000000000000000000000000000000000000000b00101600000000000000000000000000000000000000000b009e0d00000000000000000000000000000000000000000b00a71500000000000000000000000000000000000000000b00d33e00000000000000000000000000000000000000000b00851d00000000000000000000000000000000000000000b007c4000000000000000000000000000000000000000000b002f3000000000000000000000000000000000000000000b00601900000000000000000000000000000000000000000b00e13e00000000000000000000000000000000000000000b00193f00000000000000000000000000000000000000000b00ef4a00000000000000000000000000000000000000000b00021e00000000000000000000000000000000000000000b00991000000000000000000000000000000000000000000b00ce4100000000000000000000000000000000000000000b00a12f00000000000000000000000000000000000000000b00dd2b00000000000000000000000000000000000000000b005b4600000000000000000000000000000000000000000b00851300000000000000000000000000000000000000000b00522500000000000000000000000000000000000000000b008b3f00000000000000000000000000000000000000000b00d24200000000000000000000000000000000000000000b00673900000000000000000000000000000000000000000b00f60000000000000000000000000000000000000000000b00ec0800000000000000000000000000000000000000000b00dd0f00000000000000000000000000000000000000000b00cd1100000000000000000000000000000000000000000b00d31100000000000000000000000000000000000000000b00912900000000000000000000000000000000000000000b00d63c00000000000000000000000000000000000000000b00670d00000000000000000000000000000000000000000b00a54300000000000000000000000000000000000000000b00dd1100000000000000000000000000000000000000000b00334a00000000000000000000000000000000000000000b00843100000000000000000000000000000000000000000b00883100000000000000000000000000000000000000000b00cd1e00000000000000000000000000000000000000000b00b54d00000000000000000000000000000000000000000b00704600000000000000000000000000000000000000000b00ea2000000000000000000000000000000000000000000b00ae4d00000000000000000000000000000000000000000b002b0800000000000000000000000000000000000000000b00c51300000000000000000000000000000000000000000b000c0000000000000000000000000000000000000000000b00da4800000000000000000000000000000000000000000b00cc1700000000000000000000000000000000000000000b00590000000000000000000000000000000000000000000b00bd1c00000000000000000000000000000000000000000b00630600000000000000000000000000000000000000000b00a92700000000000000000000000000000000000000000b00931400000000000000000000000000000000000000000b00fa2300000000000000000000000000000000000000000b00df0800000000000000000000000000000000000000000b000e4900000000000000000000000000000000000000000b00982200000000000000000000000000000000000000000b00474a00000000000000000000000000000000000000000b00a92200000000000000000000000000000000000000000b00080000000000000000000000000000000000000000000b00280b00000000000000000000000000000000000000000b00b31b00000000000000000000000000000000000000000b004a0f00000000000000000000000000000000000000000b00644600000000000000000000000000000000000000000b008c2000000000000000000000000000000000000000000b002b0900000000000000000000000000000000000000000b00cc1a00000000000000000000000000000000000000000b00f54000000000000000000000000000000000000000000b004a1400000000000000000000000000000000000000000b00512c00000000000000000000000000000000000000000b00d20100000000000000000000000000000000000000000b00254c00000000000000000000000000000000000000000b00be4d00000000000000000000000000000000000000000b001f0100000000000000000000000000000000000000000b00011c00000000000000000000000000000000000000000b00e23200000000000000000000000000000000000000000b003e2800000000000000000000000000000000000000000b00620c00000000000000000000000000000000000000000b00304500000000000000000000000000000000000000000b000f2e00000000000000000000000000000000000000000b00f03200000000000000000000000000000000000000000b00680b00000000000000000000000000000000000000000b00904000000000000000000000000000000000000000000b00ca3f00000000000000000000000000000000000000000b00e62b00000000000000000000000000000000000000000b00ae3900000000000000000000000000000000000000000b00ff0f00000000000000000000000000000000000000000b00252c00000000000000000000000000000000000000000b003e2300000000000000000000000000000000000000000b00802300000000000000000000000000000000000000000b00293900000000000000000000000000000000000000000b00cf3600000000000000000000000000000000000000000b00e72900000000000000000000000000000000000000000b00504a00000000000000000000000000000000000000000b00a80d00000000000000000000000000000000000000000b00352c00000000000000000000000000000000000000000b00d53600000000000000000000000000000000000000000b00113700000000000000000000000000000000000000000b000a0400000000000000000000000000000000000000000b006c4000000000000000000000000000000000000000000b00933300000000000000000000000000000000000000000b00240100000000000000000000000000000000000000000b00ab0500000000000000000000000000000000000000000b00da4a00000000000000000000000000000000000000000b00b24e00000000000000000000000000000000000000000b00e24a00000000000000000000000000000000000000000b008c2800000000000000000000000000000000000000000b00912e00000000000000000000000000000000000000000b00123500000000000000000000000000000000000000000b00e34800000000000000000000000000000000000000000b00a23d00000000000000000000000000000000000000000b00de1b00000000000000000000000000000000000000000b008f3400000000000000000000000000000000000000000b007e0f00000000000000000000000000000000000000000b00a92d00000000000000000000000000000000000000000b00911500000000000000000000000000000000000000000b00804700000000000000000000000000000000000000000b007e4a00000000000000000000000000000000000000000b00a20d00000000000000000000000000000000000000000b00ec0000000000000000000000000000000000000000000b00671a00000000000000000000000000000000000000000b00cc3600000000000000000000000000000000000000000b00b12400000000000000000000000000000000000000000b000f3c00000000000000000000000000000000000000000b005b2b00000000000000000000000000000000000000000b00584700000000000000000000000000000000000000000b001d3200000000000000000000000000000000000000000b00573a00000000000000000000000000000000000000000b00e74c00000000000000000000000000000000000000000b00462c00000000000000000000000000000000000000000b007e0900000000000000000000000000000000000000000b00e50800000000000000000000000000000000000000000b008c3300000000000000000000000000000000000000000b00a00f00000000000000000000000000000000000000000b009c0500000000000000000000000000000000000000000b00c64600000000000000000000000000000000000000000b00cb3d00000000000000000000000000000000000000000b00ba0300000000000000000000000000000000000000000b00584400000000000000000000000000000000000000000b00f60600000000000000000000000000000000000000000b00a70e00000000000000000000000000000000000000000b00514200000000000000000000000000000000000000000b00a73c00000000000000000000000000000000000000000b00e32f00000000000000000000000000000000000000000b00714a00000000000000000000000000000000000000000b00e14900000000000000000000000000000000000000000b00114f00000000000000000000000000000000000000000b002c1b00000000000000000000000000000000000000000b00e32700000000000000000000000000000000000000000b00184800000000000000000000000000000000000000000b00083500000000000000000000000000000000000000000b00c20200000000000000000000000000000000000000000b00211500000000000000000000000000000000000000000b00180500000000000000000000000000000000000000000b00441300000000000000000000000000000000000000000b00294b00000000000000000000000000000000000000000b001d3500000000000000000000000000000000000000000b00081a00000000000000000000000000000000000000000b00320700000000000000000000000000000000000000000b006e3a00000000000000000000000000000000000000000b00740700000000000000000000000000000000000000000b00263f00000000000000000000000000000000000000000b002d3300000000000000000000000000000000000000000b00e14100000000000000000000000000000000000000000b000d0a00000000000000000000000000000000000000000b00382800000000000000000000000000000000000000000b00481900000000000000000000000000000000000000000b00312400000000000000000000000000000000000000000b00b62d00000000000000000000000000000000000000000b00541100000000000000000000000000000000000000000a00f00f00000000000000000000000000000000000000000a00201000000000000000000000000000000000000000000a00501000000000000000000000000000000000000000000b00f10600000000000000000000000000000000000000000b00ef3700000000000000000000000000000000000000000b00082f00000000000000000000000000000000000000000b00911900000000000000000000000000000000000000000b009a1900000000000000000000000000000000000000000b003b2f00000000000000000000000000000000000000000b00991600000000000000000000000000000000000000000b00cb4700000000000000000000000000000000000000000300326501000000000000000000000000000000000000000300a0a201000000000000000000000000000000000000000300aea201000000000000000000000000000000000000000300b0a201000000000000000000000000000000000000000300f2a301000000000000000000000000000000000000000300d6a5010000000000000000000000000000000000000003002ca601000000000000000000000000000000000000000300a4a901000000000000000000000000000000000000000300b2a90100000000000000000000000000000000000000030030ab0100000000000000000000000000000000000000030042ab0100000000000000000000000000000000000000030054ab0100000000000000000000000000000000000000030062ab0100000000000000000000000000000000000000030070ab01000000000000000000000000000000000000000300e0ab010000000000000000000000000000000000000003009cad0100000000000000000000000000000000000000030050ae0100000000000000000000000000000000000000030088ae0100000000000000000000000000000000000000030092ae0100000000000000000000000000000000000000030048af0100000000000000000000000000000000000000030082af01000000000000000000000000000000000000000300a2b001000000000000000000000000000000000000000300a2b1010000000000000000000000000000000000000003003ab20100000000000000000000000000000000000000030048b201000000000000000000000000000000000000000300bab2010000000000000000000000000000000000000003002cb30100000000000000000000000000000000000000030042b301000000000000000000000000000000000000000300e4b30100000000000000000000000000000000000000030054b401000000000000000000000000005e6500000400f1ff000000000000000000000000000000006465000000000300268302000000000000000000000000006765000000000300f48302000000000000000000000000006a650000000003001c8802000000000000000000000000006d65000000000300428802000000000000000000000000007065000000000300f28302000000000000000000000000007465000000000300e28302000000000000000000000000007865000000000300188802000000000000000000000000007d65000000000300d08402000000000000000000000000008265000000000300188402000000000000000000000000008765000000000300ba8602000000000000000000000000008c65000000000300148402000000000000000000000000009165000000000300e48402000000000000000000000000009665000000000300908402000000000000000000000000009b650000000003004e840200000000000000000000000000a06500000000030052870200000000000000000000000000a5650000000003005e840200000000000000000000000000aa65000000000300b6840200000000000000000000000000af65000000000300c2840200000000000000000000000000b465000000000300a4860200000000000000000000000000b96500000000030098850200000000000000000000000000be6500000000030082870200000000000000000000000000c365000000000300c4860200000000000000000000000000c8650000000003002e850200000000000000000000000000cd6500000000030032860200000000000000000000000000d2650000000003007a860200000000000000000000000000d765000000000300a0860200000000000000000000000000dc65000000000300c6840200000000000000000000000000e165000000000300e6860200000000000000000000000000e6650000000003005c870200000000000000000000000000eb65000000000300ac870200000000000000000000000000f0650000000003002c840200000000000000000000000000f56500000000030032880200000000000000000000000000fb650000000003003688020000000000000000000000000001660000000003001e8802000000000000000000000000000766000000000300228902000000000000000000000000000d66000000000300028a020000000000000000000000000013660000000003002689020000000000000000000000000019660000000003008e8902000000000000000000000000001f66000000000300088a02000000000000000000000000002566000000000300048a02000000000000000000000000002b66000000000300a488020000000000000000000000000031660000000003007889020000000000000000000000000037660000000003001e8a02000000000000000000000000003d660000000003004489020000000000000000000000000043660000000003003e89020000000000000000000000000049660000000003000e8a02000000000000000000000000004f66000000000300628902000000000000000000000000005566000000000300228a02000000000000000000000000005b66000000000300a68902000000000000000000000000006166000000000300a08902000000000000000000000000006766000000000300128a02000000000000000000000000006d66000000000300ce8902000000000000000000000000007366000000000300f08902000000000000000000000000007966000000000300ee8902000000000000000000000000007f66000000000300ea8902000000000000000000000000008566000000000300588902000000000000000000000000008b66000000000300b8890200000000000000000000000000a7660000020203004288020000000000e601000000000000af66000002020300f4830200000000002804000000000000b6660000020203001c880200000000002600000000000000bd660000020203002683020000000000ce000000000000009166000012000300c845010000000000861e000000000000a066000010000300cc340100000000000000000000000000002e726f64617461002e65685f6672616d65002e74657874002e7364617461002e64617461002e627373002e64656275675f616262726576002e64656275675f696e666f002e64656275675f6172616e676573002e64656275675f72616e676573002e64656275675f737472002e64656275675f7075626e616d6573002e64656275675f7075627479706573002e72697363762e61747472696275746573002e64656275675f6c696e65002e636f6d6d656e74002e73796d746162002e7368737472746162002e73747274616200007374616b655f736d742e386464326133386433633037646163632d6367752e30002e4c435049305f30005f5a4e34636f72653370747231373364726f705f696e5f706c616365244c5424616c6c6f632e2e7665632e2e696e746f5f697465722e2e496e746f49746572244c5424244c502424753562247538247533622424753230243230247535642424432424753562247538247533622424753230243332247535642424432461786f6e5f74797065732e2e67656e6572617465642e2e7374616b655f7265616465722e2e5374616b65496e666f44656c74612452502424475424244754243137683437613765613563366266363330356645002e4c706372656c5f686930005f5a4e36345f244c5424616c6c6f632e2e72632e2e5263244c54245424475424247532302461732475323024636f72652e2e6f70732e2e64726f702e2e44726f70244754243464726f703137683663346239333364656266363135663545005f5f727573745f6465616c6c6f63005f5a4e34636f726533707472343664726f705f696e5f706c616365244c5424616c6c6f632e2e7665632e2e566563244c5424753824475424244754243137683635613963343931333965643939373745005f5a4e34636f726533707472383864726f705f696e5f706c616365244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e7365742e2e4254726565536574244c54247574696c2e2e736d742e2e4c6f636b496e666f24475424244754243137683438613635376438646464366532326245002e4c706372656c5f686931002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e30005f5a4e34636f72653970616e69636b696e673570616e69633137686437373538656430613265383739363145005f5a4e35616c6c6f633131636f6c6c656374696f6e733562747265653373657432314254726565536574244c542454244324412447542436696e736572743137683132343337323662373533323537373145005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565367365617263683134325f244c5424696d706c2475323024616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e4e6f6465526566244c5424426f72726f77547970652443244b24432456244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4c6561664f72496e7465726e616c244754242447542431317365617263685f747265653137683331653862613736663538633563313145005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f646532314c6561664e6f6465244c54244b2443245624475424336e65773137683339666330303661613430353065373245005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f64653235496e7465726e616c4e6f6465244c54244b2443245624475424336e65773137683731366362643563613232623662316645005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f646532313448616e646c65244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e4e6f6465526566244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4d75742443244b24432456244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e496e7465726e616c24475424244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e45646765244754243130696e736572745f6669743137686133363335336433636163353566646545002e4c706372656c5f686934002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e3639002e4c706372656c5f686935002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e3635005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243135636f70795f66726f6d5f736c69636531376c656e5f6d69736d617463685f6661696c3137686531663934356265353831313135613845002e4c706372656c5f686936002e4c706372656c5f686932002e4c706372656c5f686933002e4c706372656c5f686937002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e3537002e4c706372656c5f686938005f5f727573745f616c6c6f63005f5f727573745f616c6c6f635f6572726f725f68616e646c6572005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b2443245624475424313562756c6b5f737465616c5f6c6566743137683831346639376465613163366363333245002e4c706372656c5f686939002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e3733002e4c706372656c5f68693131002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e3735002e4c706372656c5f68693130002e4c706372656c5f68693132002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e3737005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b2443245624475424313662756c6b5f737465616c5f72696768743137686563303938393134323636343965323345002e4c706372656c5f68693133002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e3830002e4c706372656c5f68693135002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e3832002e4c706372656c5f68693134002e4c706372656c5f68693136005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b244324562447542432356d657267655f747261636b696e675f6368696c645f656467653137683962653866643964663537626138333045002e4c706372656c5f68693138002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e3835002e4c706372656c5f68693137002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e3837005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b244324562447542438646f5f6d657267653137683766313436336161373166393732393645002e4c706372656c5f68693139005f5a4e35616c6c6f633131636f6c6c656374696f6e733562747265653672656d6f76653235395f244c5424696d706c2475323024616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e48616e646c65244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e4e6f6465526566244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4d75742443244b24432456244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4c65616624475424244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4b562447542424475424313472656d6f76655f6c6561665f6b763137683430313336343539653762343932393945005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f64653132354e6f6465526566244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4d75742443244b24432456244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4c6561664f72496e7465726e616c24475424313663686f6f73655f706172656e745f6b763137683664396533663635623666653665643145002e4c706372656c5f68693230005f5a4e37636b625f73746433656e7634415247563137683861626337373932303633656163623745005f5a4e35616c6c6f63377261775f7665633139526177566563244c54245424432441244754243131616c6c6f636174655f696e3137683961373435623837316432623838663945002e4c706372656c5f68693231002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e383436002e4c706372656c5f68693233002e4c706372656c5f68693232002e4c424231335f3138002e4c706372656c5f68693234002e4c706372656c5f68693235002e4c706372656c5f68693236005f5a4e34636f726535736c69636535696e64657837345f244c5424696d706c2475323024636f72652e2e6f70732e2e696e6465782e2e496e646578244c542449244754242475323024666f72247532302424753562245424753564242447542435696e6465783137683064326565363561653136626361336545005f5a4e3131315f244c5424616c6c6f632e2e7665632e2e566563244c54245424475424247532302461732475323024616c6c6f632e2e7665632e2e737065635f66726f6d5f697465725f6e65737465642e2e5370656346726f6d497465724e6573746564244c5424542443244924475424244754243966726f6d5f697465723137683032353562336632346332623633633445005f5a4e35616c6c6f63337665633136566563244c542454244324412447542434707573683137683832346530366138613965323339383745005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f7233616e793137683031323866356465313834336464653445002e4c706372656c5f68693238002e4c706372656c5f68693237005f5a4e3130325f244c5424636b625f7374616e64616c6f6e655f74797065732e2e67656e6572617465642e2e626c6f636b636861696e2e2e42797465735265616465722475323024617324753230246d6f6c6563756c652e2e7072656c7564652e2e52656164657224475424367665726966793137683135663233383466353032373265326345005f5a4e386d6f6c6563756c6535627974657335427974657335736c6963653137683133633337653065643765643238336345005f5a4e3230636b625f7374616e64616c6f6e655f74797065733967656e6572617465643130626c6f636b636861696e354279746573387261775f646174613137686165613062386538653731396665363945005f5a4e37636b625f7374643130686967685f6c6576656c31396c6f61645f63656c6c5f747970655f686173683137683563643636373336663632346636613545002e4c706372656c5f68693330002e4c4a544931335f30002e4c424231335f3732005f5a4e347574696c3668656c70657231386765745f7374616b655f736d745f646174613137683066643534393634653339306137323245005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231365374616b65536d7443656c6c4461746131366d657461646174615f747970655f69643137683333316537333761333766666465306145005f5a4e347574696c3668656c70657232366765745f6d65746164615f646174615f62795f747970655f69643137686130366330323062366338343062303345005f5a4e396d6f6c6563756c65323672656164657236437572736f72323164796e7665635f736c6963655f62795f696e6465783137683464633230383535323662653634303045005f5a4e347574696c3668656c70657232376765745f63656c6c5f636f756e745f62795f747970655f686173683137683433316433366633633236643131663045002e4c424231335f3933002e4c424231335f3934005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f72656164657237547970654964733134787564745f747970655f686173683137686334653636633566343738343237356145005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f726561646572375479706549647331397374616b655f736d745f636f64655f686173683137683939313230643232643561376161363745005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f726561646572375479706549647331377374616b655f736d745f747970655f69643137683133613730383736373561386135323245005f5a4e347574696c3668656c70657231356765745f7363726970745f686173683137686133663334636563626161396538326445005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f72656164657237547970654964733230636865636b706f696e745f636f64655f686173683137683561366363373337366465333564383045005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f72656164657237547970654964733138636865636b706f696e745f747970655f69643137683062376537323033303666383865346345005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f7265616465723754797065496473313877697468647261775f636f64655f686173683137686636356461336666633664366137323445005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f726561646572375479706549647331386d657461646174615f636f64655f686173683137683263623137613437626166656264306645005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f726561646572375479706549647331366d657461646174615f747970655f69643137683833306539326563613930383864363745005f5a4e3230636b625f7374616e64616c6f6e655f74797065733967656e6572617465643130626c6f636b636861696e31315769746e65737341726773346c6f636b3137686233326333343036613431316531636245005f5a4e39385f244c54246d6f6c6563756c65322e2e7265616465722e2e437572736f72247532302461732475323024636f72652e2e636f6e766572742e2e46726f6d244c5424616c6c6f632e2e7665632e2e566563244c542475382447542424475424244754243466726f6d3137686365383937663564613837343036643045005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231345374616b65496e666f44656c7461313169735f696e6372656173653137683166386136356661303836623163316645005f5a4e347574696c3668656c70657231376765745f63757272656e745f65706f63683137683561353332396138346166353437623445005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231385374616b65536d74557064617465496e666f3135616c6c5f7374616b655f696e666f733137686331656532343334363962343463366245005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231305374616b65496e666f73336c656e3137683862303137666338646362303233393945005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231305374616b65496e666f73336765743137683536663765343736643831623335613045005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f726561646572395374616b65496e666f34616464723137683737663935343236353164653934373045005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231345374616b65496e666f44656c746136616d6f756e743137683736303137613463316430633135626445005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231385374616b65536d74557064617465496e666f31356f6c645f65706f63685f70726f6f663137683835396638343561623737663561346545005f5a4e347574696c33736d7431317536345f746f5f683235363137686135386530356361383833323362356245005f5a4e347574696c33736d7431377665726966795f326c617965725f736d743137683530613034653963613062323634646445005f5a4e347574696c3668656c70657232326765745f7374616b655f7570646174655f696e666f733137686566336433396666393563396264616445005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231345374616b65496e666f44656c74613138696e61756775726174696f6e5f65706f63683137683538323561303933383837366165313345005f5a4e347574696c3668656c70657233306765745f7374616b655f61745f646174615f62795f6c6f636b5f686173683137686361666239343538306137663634303645005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231355374616b65417443656c6c446174613564656c74613137683762333332613765343438316530613845005f5a4e3130385f244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6d61702e2e49746572244c54244b2443245624475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683436323362663162343430666237623945005f5a4e347574696c3668656c706572323563616c635f7769746864726177616c5f6c6f636b5f686173683137686337616539656536383134393866383145005f5a4e347574696c3668656c70657233336765745f77697468647261775f61745f646174615f62795f6c6f636b5f686173683137683632306461356439643938323335613245005f5a4e347574696c3668656c70657231356765745f71756f72756d5f73697a653137686634656138393232363736633436333645005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231385374616b65536d74557064617465496e666f31356e65775f65706f63685f70726f6f663137686236623761343265306435646564653745002e4c706372656c5f68693239002e4c706372656c5f68693433007374722e31002e4c424231335f323739005f5a4e34636f72653970616e69636b696e673970616e69635f666d743137686436616161656662346334646538633945002e4c706372656c5f68693331002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e3436002e4c706372656c5f68693332002e4c616e6f6e2e63396664323635383763663061663763663065366537386464383734316533382e33002e4c706372656c5f68693333002e4c706372656c5f68693334002e4c616e6f6e2e30656130363565396135373639326336653434396165616266643062303633332e3139005f5a4e34636f726536726573756c743133756e777261705f6661696c65643137683030653934303161326339653536633045002e4c706372656c5f68693435002e4c706372656c5f68693436002e4c706372656c5f68693335002e4c706372656c5f68693336002e4c616e6f6e2e63396664323635383763663061663763663065366537386464383734316533382e34002e4c706372656c5f68693337002e4c706372656c5f68693338002e4c706372656c5f68693339002e4c706372656c5f68693430002e4c706372656c5f68693431002e4c706372656c5f68693432002e4c706372656c5f68693434002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e363300727573745f626567696e5f756e77696e64005f5a4e37636b625f7374643873797363616c6c73366e617469766534657869743137686334346330613764356530656238316345005f5a4e397374616b655f736d7431316f6f6d5f68616e646c65723137686333633466356639346562636164656245005f5f72675f6f6f6d005f5f72675f616c6c6f63005f5a4e3130365f244c542462756464795f616c6c6f632e2e6e6f6e5f746872656164736166655f616c6c6f632e2e4e6f6e54687265616473616665416c6c6f63247532302461732475323024636f72652e2e616c6c6f632e2e676c6f62616c2e2e476c6f62616c416c6c6f632447542435616c6c6f633137683966656332343337626566343266383945005f5f72675f6465616c6c6f63005f5a4e3130365f244c542462756464795f616c6c6f632e2e6e6f6e5f746872656164736166655f616c6c6f632e2e4e6f6e54687265616473616665416c6c6f63247532302461732475323024636f72652e2e616c6c6f632e2e676c6f62616c2e2e476c6f62616c416c6c6f6324475424376465616c6c6f633137686530336235656339643238613732396445005f5f72675f7265616c6c6f63005f5f72675f616c6c6f635f7a65726f6564005f5f727573745f7265616c6c6f63005f5f727573745f616c6c6f635f7a65726f6564005f5a4e35616c6c6f63377261775f766563313763617061636974795f6f766572666c6f773137683736396433373734353939336431626545005f5a4e396d6f6c6563756c6532367265616465723130385f244c5424696d706c2475323024636f72652e2e636f6e766572742e2e46726f6d244c54246d6f6c6563756c65322e2e7265616465722e2e437572736f72244754242475323024666f722475323024616c6c6f632e2e7665632e2e566563244c5424753824475424244754243466726f6d3137683965653331373661666261663535343545002e4c706372656c5f68693437002e4c706372656c5f68693438002e4c706372656c5f68693439002e4c706372656c5f68693530002e4c706372656c5f68693531002e4c706372656c5f68693532002e4c706372656c5f68693533002e4c706372656c5f68693534002e4c706372656c5f68693535002e4c706372656c5f68693536002e4c706372656c5f68693537002e4c706372656c5f68693538002e4c706372656c5f68693539002e4c706372656c5f68693630002e4c706372656c5f68693631002e4c706372656c5f68693632005f5a4e396d6f6c6563756c65323672656164657238355f244c5424696d706c2475323024636f72652e2e636f6e766572742e2e46726f6d244c54246d6f6c6563756c65322e2e7265616465722e2e437572736f72244754242475323024666f7224753230247538244754243466726f6d3137686461653235633931336631613435396545002e4c706372656c5f68693633002e4c706372656c5f68693634002e4c706372656c5f68693635002e4c706372656c5f68693636005f5a4e396d6f6c6563756c65323672656164657238365f244c5424696d706c2475323024636f72652e2e636f6e766572742e2e46726f6d244c54246d6f6c6563756c65322e2e7265616465722e2e437572736f72244754242475323024666f722475323024753634244754243466726f6d3137686232663035653938653831303635333145002e4c706372656c5f68693637002e4c706372656c5f68693638002e4c706372656c5f68693639002e4c706372656c5f68693730002e4c706372656c5f68693731002e4c706372656c5f68693732002e4c706372656c5f68693733002e4c706372656c5f68693734005f5a4e396d6f6c6563756c65323672656164657236437572736f723876616c69646174653137683930306131623931383065653939313845005f5a4e396d6f6c6563756c65323672656164657236437572736f7231346765745f6974656d5f636f756e743137683362393033346337303939633162346445002e4c706372656c5f68693735002e4c706372656c5f68693736002e4c706372656c5f68693737002e4c706372656c5f68693738002e4c706372656c5f68693739002e4c706372656c5f68693830005f5a4e396d6f6c6563756c65323672656164657236437572736f723139636f6e766572745f746f5f72617762797465733137683634326263616436376665326537643145002e4c706372656c5f68693831002e4c706372656c5f68693832002e4c706372656c5f68693833002e4c706372656c5f68693834002e4c706372656c5f68693835002e4c706372656c5f68693836002e4c706372656c5f68693837002e4c706372656c5f68693838005f5a4e3131626c616b6532625f72656637777261707065723134426c616b6532624275696c646572356275696c643137683964636431366662373535323133626345005f5a4e3131626c616b6532625f7265663131626c616b6532625f7265663138626c616b6532625f696e69745f706172616d3137683431613831343963666239633164343445005f5a4e3131626c616b6532625f7265663131626c616b6532625f7265663134626c616b6532625f7570646174653137683337646637643338333264666265336545002e4c706372656c5f68693839005f5a4e3131626c616b6532625f7265663131626c616b6532625f7265663130626c616b6532625f49563137686532356438333932346363316638393145005f5a4e3131626c616b6532625f7265663131626c616b6532625f7265663136626c616b6532625f636f6d70726573733137683531363361326435303733336262323945002e4c43504935315f30002e4c43504935315f31002e4c43504935315f32002e4c43504935315f33002e4c43504935315f34002e4c43504935315f35002e4c43504935315f36002e4c43504935315f37002e4c706372656c5f68693930002e4c706372656c5f68693931002e4c706372656c5f68693932002e4c706372656c5f68693933002e4c706372656c5f68693934002e4c706372656c5f68693935002e4c706372656c5f68693936002e4c706372656c5f68693937005f5a4e3131626c616b6532625f726566377772617070657237426c616b6532623866696e616c697a653137683431356365303263316365386263623745005f5a4e313162756464795f616c6c6f63313162756464795f616c6c6f6331304275646479416c6c6f63336e65773137683039343964346234353436656265666245005f5a4e313162756464795f616c6c6f63313162756464795f616c6c6f6337726f756e6475703137686533656266373734346663663366363345002e4c706372656c5f6869313035007374722e342e3631005f5a4e313162756464795f616c6c6f63313162756464795f616c6c6f63366e626c6f636b3137683537623963376462363561386133343745005f5a4e313162756464795f616c6c6f63313162756464795f616c6c6f6331304275646479416c6c6f633131626c6f636b5f696e6465783137683333633165376336333564613363643945005f5a4e34636f7265366f7074696f6e31336578706563745f6661696c65643137686332333330616533386638616564396545002e4c706372656c5f6869313130002e4c706372656c5f6869313036002e4c706372656c5f6869313037002e4c706372656c5f68693938002e4c706372656c5f6869313030007374722e322e3632002e4c706372656c5f6869313031007374722e332e3633002e4c706372656c5f6869313032002e4c706372656c5f6869313033007374722e312e3630002e4c706372656c5f6869313034002e4c706372656c5f6869313131002e4c706372656c5f6869313038007374722e302e3539002e4c706372656c5f68693939002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3135002e4c706372656c5f6869313132002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3238005f5a4e34636f72653970616e69636b696e67313370616e69635f646973706c61793137683538303536323433613031393534316645002e4c706372656c5f6869313039002e4c706372656c5f6869313133002e4c706372656c5f6869313134002e4c706372656c5f6869313135002e4c706372656c5f6869313136002e4c706372656c5f6869313137002e4c706372656c5f6869313139002e4c706372656c5f6869313230002e4c706372656c5f6869313138002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3338005f5a4e313162756464795f616c6c6f633130666173745f616c6c6f633946617374416c6c6f63336e65773137683239303962396561363461333531383845002e4c706372656c5f6869313232002e4c706372656c5f6869313231002e4c706372656c5f6869313233002e4c706372656c5f6869313234005f5a4e397374616b655f736d7435414c4c4f433137686638616535353638343561346431386345002e4c706372656c5f6869313238002e4c706372656c5f6869313333002e4c706372656c5f6869313334002e4c706372656c5f6869313331002e4c706372656c5f6869313335002e4c706372656c5f6869313336002e4c706372656c5f6869313332002e4c706372656c5f6869313237002e4c706372656c5f6869313239002e4c706372656c5f6869313330002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e32002e4c706372656c5f6869313235002e4c706372656c5f6869313236002e4c706372656c5f6869313337002e4c706372656c5f6869313338002e4c706372656c5f6869313339002e4c706372656c5f6869313433002e4c706372656c5f6869313432002e4c706372656c5f6869313436002e4c706372656c5f6869313438002e4c706372656c5f6869313439002e4c706372656c5f6869313530002e4c706372656c5f6869313437002e4c706372656c5f6869313430002e4c706372656c5f6869313431002e4c706372656c5f6869313434002e4c706372656c5f6869313435005f5a4e35616c6c6f63377261775f7665633139526177566563244c54245424432441244754243131616c6c6f636174655f696e3137683334393639363464643031633234363645005f5a4e35616c6c6f63377261775f7665633139526177566563244c542454244324412447542437726573657276653231646f5f726573657276655f616e645f68616e646c653137686234636364626536643135363830353445002e4c706372656c5f6869313531007374722e302e3639005f5a4e35616c6c6f63377261775f7665633139526177566563244c5424542443244124475424313467726f775f616d6f7274697a65643137683131313435313531653037646531613245005f5a4e35616c6c6f63377261775f766563313166696e6973685f67726f773137683362363537323731663362336132663345005f5a4e35616c6c6f63377261775f7665633139526177566563244c54245424432441244754243136726573657276655f666f725f707573683137683364383734353931323332303230376445002e4c706372656c5f6869313532002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e313734002e4c706372656c5f6869313533002e4c706372656c5f6869313534005f5a4e3230636b625f7374616e64616c6f6e655f74797065733130636f6e76657273696f6e3130626c6f636b636861696e3134395f244c5424696d706c2475323024636b625f7374616e64616c6f6e655f74797065732e2e7072656c7564652e2e5061636b244c5424636b625f7374616e64616c6f6e655f74797065732e2e67656e6572617465642e2e626c6f636b636861696e2e2e427974653332244754242475323024666f72247532302424753562247538247533622424753230243332247535642424475424347061636b3137683838633365666265633136666335636345005f5a4e3230636b625f7374616e64616c6f6e655f74797065733130636f6e76657273696f6e397072696d69746976653133365f244c5424696d706c2475323024636b625f7374616e64616c6f6e655f74797065732e2e7072656c7564652e2e5061636b244c5424636b625f7374616e64616c6f6e655f74797065732e2e67656e6572617465642e2e626c6f636b636861696e2e2e4279746573244754242475323024666f72247532302424753562247538247535642424475424347061636b3137686534363231633861323935306563356145005f5a4e3133325f244c5424616c6c6f632e2e7665632e2e566563244c5424542443244124475424247532302461732475323024616c6c6f632e2e7665632e2e737065635f657874656e642e2e53706563457874656e64244c54242452462454244324636f72652e2e736c6963652e2e697465722e2e49746572244c5424542447542424475424244754243131737065635f657874656e643137683464663561353366366631653763336445002e4c706372656c5f6869313535007374722e322e3638005f5a4e39375f244c5424636b625f7374616e64616c6f6e655f74797065732e2e67656e6572617465642e2e626c6f636b636861696e2e2e5363726970742475323024617324753230246d6f6c6563756c652e2e7072656c7564652e2e456e746974792447542431316e65775f6275696c6465723137683663323863633439326130386634363645005f5a4e3130355f244c5424636b625f7374616e64616c6f6e655f74797065732e2e67656e6572617465642e2e626c6f636b636861696e2e2e5363726970744275696c6465722475323024617324753230246d6f6c6563756c652e2e7072656c7564652e2e4275696c64657224475424356275696c643137683462313334356436646334623638326145002e4c706372656c5f6869313536002e4c706372656c5f6869313537002e4c706372656c5f6869313538005f5a4e36315f244c5424636b625f7374642e2e6572726f722e2e5379734572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137686534313062343262643137646531353845002e4c706372656c5f6869313539002e4c4a544937375f30002e4c424237375f31002e4c706372656c5f6869313630002e4c616e6f6e2e35366333623930656239393266643662383361623665306438306633656532622e3339002e4c424237375f32002e4c706372656c5f6869313631002e4c616e6f6e2e35366333623930656239393266643662383361623665306438306633656532622e3338002e4c424237375f33002e4c706372656c5f6869313632002e4c616e6f6e2e35366333623930656239393266643662383361623665306438306633656532622e3336002e4c706372656c5f6869313633002e4c616e6f6e2e35366333623930656239393266643662383361623665306438306633656532622e3337002e4c424237375f34002e4c706372656c5f6869313634002e4c424237375f36002e4c706372656c5f6869313635002e4c616e6f6e2e35366333623930656239393266643662383361623665306438306633656532622e3333002e4c706372656c5f6869313636002e4c616e6f6e2e35366333623930656239393266643662383361623665306438306633656532622e3334005f5a4e34636f726533666d7439466f726d6174746572323564656275675f7475706c655f6669656c64315f66696e6973683137683963326264643732306464613133376545005f5a4e34636f726533707472323864726f705f696e5f706c616365244c542424524624753634244754243137683135383466626334313265393865303445005f5a4e37636b625f7374643130686967685f6c6576656c31396c6f61645f63656c6c5f6c6f636b5f686173683137683339633636646239366138646337393445005f5a4e37636b625f7374643130686967685f6c6576656c31346c6f61645f63656c6c5f646174613137683061353964663134343334336539316145005f5a4e34636f7265336f70733866756e6374696f6e36466e4f6e63653963616c6c5f6f6e63653137683331326365396462383432326365623645005f5a4e34636f72653370747231303264726f705f696e5f706c616365244c542424524624636f72652e2e697465722e2e61646170746572732e2e636f706965642e2e436f70696564244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c542475382447542424475424244754243137683465633534623435323134663763393045002e4c43504938365f30005f5a4e34636f726533666d74336e756d33696d7037666d745f7536343137683238366534643532373433386334363745002e4c706372656c5f6869313637002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333234002e4c706372656c5f6869313638002e4c706372656c5f6869313639002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e3233005f5a4e34636f726533666d7439466f726d617474657231327061645f696e74656772616c3137686238656639343965396131613633346545005f5a4e34636f726533666d7439466f726d617474657231327061645f696e74656772616c313277726974655f7072656669783137683834663538656430383761336264393345002e4c43504938395f30002e4c43504938395f31005f5a4e34636f726533666d7439466f726d6174746572337061643137683433336537613934646232626438653245002e4c706372656c5f6869313730002e4c706372656c5f6869313731005f5a4e34636f726533666d743577726974653137683537653362636463656237646630393145002e4c706372656c5f6869313732005f5a4e36305f244c5424636f72652e2e63656c6c2e2e426f72726f774572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137686163386261333334363731373261333845002e4c706372656c5f6869313733002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e313730005f5a4e36335f244c5424636f72652e2e63656c6c2e2e426f72726f774d75744572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683636336332373865383138373636393045002e4c706372656c5f6869313734002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e313731005f5a4e34636f726533666d74336e756d35335f244c5424696d706c2475323024636f72652e2e666d742e2e4c6f7765724865782475323024666f7224753230246936342447542433666d743137686632356530653835343735353364373145002e4c706372656c5f6869313735002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333232002e4c43504939375f30002e4c43504939375f31002e4c43504939375f32005f5a4e36385f244c5424636f72652e2e666d742e2e6275696c646572732e2e50616441646170746572247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f7374723137686539366438303337316562386433343445002e4c706372656c5f6869313736002e4c706372656c5f6869313737002e4c706372656c5f6869313738002e4c706372656c5f6869313739005f5a4e34636f726533666d74355772697465313077726974655f636861723137686664666234386663643336373461323845005f5a4e34636f726533666d743557726974653977726974655f666d743137683364623431343565346436363932376245002e4c706372656c5f6869313830002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333237005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f7374723137683865303931326361326264646233386345005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e577269746524475424313077726974655f636861723137683239666437616639333939643762333645005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f666d743137683565373464633863623261616161323645002e4c706372656c5f6869313831005f5a4e34636f726533666d74386275696c64657273313044656275675475706c65356669656c643137686134393061356537663734366534656245002e4c706372656c5f6869313833002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e323933002e4c706372656c5f6869313834002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333030002e4c706372656c5f6869313832002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333031002e4c706372656c5f6869313835002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e323839002e4c706372656c5f6869313836002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e323932005f5a4e34636f726533666d74386275696c6465727338446562756753657435656e7472793137686531623638303262326163636539656445002e4c706372656c5f6869313930002e4c706372656c5f6869313838002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333033002e4c706372656c5f6869313837002e4c706372656c5f6869313839002e4c706372656c5f6869313932002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333032002e4c706372656c5f6869313931002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e313537005f5a4e34636f726533666d74336e756d35325f244c5424696d706c2475323024636f72652e2e666d742e2e55707065724865782475323024666f72247532302469382447542433666d743137683438643832613435336137306166353745002e4c706372656c5f6869313933005f5a4e34636f726533666d74336e756d35325f244c5424696d706c2475323024636f72652e2e666d742e2e4c6f7765724865782475323024666f72247532302469382447542433666d743137683039663834613031663936303437366145002e4c706372656c5f6869313934005f5a4e34325f244c54242452462454247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137686332303631326561373836393861653445002e4c706372656c5f6869313935002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333337005f5a4e36375f244c5424636f72652e2e61727261792e2e54727946726f6d536c6963654572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683532646436363362353834636335356645002e4c706372656c5f6869313936002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e353537002e4c706372656c5f6869313937002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e353333002e4c706372656c5f6869313939002e4c706372656c5f6869313938005f5a4e34636f726533666d74336e756d35335f244c5424696d706c2475323024636f72652e2e666d742e2e55707065724865782475323024666f7224753230246936342447542433666d743137683464336136353331313038303933376445002e4c706372656c5f6869323030005f5a4e35616c6c6f63377261775f7665633139526177566563244c542454244324412447542437726573657276653231646f5f726573657276655f616e645f68616e646c653137686332663335393562613638613033633645005f5a4e34325f244c54242452462454247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683035646461313430303562373034353645005f5a4e34325f244c54242452462454247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683431323134373832613466363464656645005f5a4e36355f244c5424616c6c6f632e2e7665632e2e566563244c5424542443244124475424247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137686464613861616433336135376363313045002e4c706372656c5f6869323031002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e323533002e4c706372656c5f6869323032002e4c706372656c5f6869323033002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333038005f5a4e35616c6c6f63337665633136566563244c54245424432441244754243131657874656e645f776974683137683935323361376565386561616133316645005f5a4e35616c6c6f63377261775f7665633139526177566563244c542454244324412447542437726573657276653231646f5f726573657276655f616e645f68616e646c653137686534386235666233366361343936633545005f5a4e35616c6c6f63377261775f766563313166696e6973685f67726f773137686465323762646133633136313431313345005f5a4e396d6f6c6563756c65323672656164657237726561645f61743137686436323832346538376630396538383045002e4c706372656c5f6869323133007374722e312e333034002e4c706372656c5f6869323036002e4c706372656c5f6869323037002e4c706372656c5f6869323034002e4c706372656c5f6869323035002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e31002e4c706372656c5f6869323132002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3136002e4c706372656c5f6869323134002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3139002e4c706372656c5f6869323038002e4c706372656c5f6869323039002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e36002e4c706372656c5f6869323130002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3132002e4c706372656c5f6869323131002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3134005f5a4e36315f244c54246d6f6c6563756c65322e2e7265616465722e2e4572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683238346238363235356264316239336545002e4c706372656c5f6869323135002e4c7377697463682e7461626c652e5f5a4e36315f244c54246d6f6c6563756c65322e2e7265616465722e2e4572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683238346238363235356264316239336545002e4c706372656c5f6869323136002e4c7377697463682e7461626c652e5f5a4e36315f244c54246d6f6c6563756c65322e2e7265616465722e2e4572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d7431376832383462383632353562643162393365452e343137002e4c706372656c5f6869323139002e4c706372656c5f6869323137002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e32002e4c706372656c5f6869323138002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e33002e4c706372656c5f6869323230002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3238005f5a4e396d6f6c6563756c65323672656164657236437572736f723133756e7061636b5f6e756d6265723137683635326430373132666263326536343145002e4c706372656c5f6869323231002e4c706372656c5f6869323232002e4c706372656c5f6869323233002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3331002e4c706372656c5f6869323234002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3335002e4c706372656c5f6869323331002e4c706372656c5f6869323235002e4c706372656c5f6869323236002e4c706372656c5f6869323330002e4c706372656c5f6869323237002e4c706372656c5f6869323238002e4c706372656c5f6869323239002e4c706372656c5f6869323332002e4c706372656c5f6869323333002e4c706372656c5f6869323334002e4c706372656c5f6869323335002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3430002e4c706372656c5f6869323336002e4c706372656c5f6869323337002e4c706372656c5f6869323338002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3538002e4c706372656c5f6869323339002e4c706372656c5f6869323430002e4c706372656c5f6869323431002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3634005f5a4e36395f244c5424616c6c6f632e2e7665632e2e566563244c54247538244754242475323024617324753230246d6f6c6563756c65322e2e7265616465722e2e526561642447542434726561643137683538323363346134366134643066373445002e4c706372656c5f6869323432002e4c706372656c5f6869323433002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3638005f5a4e34636f726533707472343664726f705f696e5f706c616365244c5424616c6c6f632e2e7665632e2e566563244c5424753824475424244754243137683139303635656264313265376238616645005f5a4e31387370617273655f6d65726b6c655f74726565346832353634483235363131706172656e745f706174683137683635373836666235326663646564306445005f5a4e37305f244c54247370617273655f6d65726b6c655f747265652e2e747265652e2e4272616e63684b6579247532302461732475323024636f72652e2e636d702e2e4f72642447542433636d703137683263653439633663323334323262346545005f5a4e39385f244c5424636b625f7374642e2e686967685f6c6576656c2e2e517565727949746572244c54244624475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683764366161393561356131323831396645002e4c706372656c5f6869323434007374722e302e333431002e4c706372656c5f6869323436002e4c706372656c5f6869323435005f5a4e35616c6c6f6335626f7865643136426f78244c542454244324412447542431336e65775f756e696e69745f696e3137683364666539356665666465623631663145005f5a4e35616c6c6f6335626f7865643136426f78244c542454244324412447542431336e65775f756e696e69745f696e3137683664383831353535333436643564303245005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f646532313448616e646c65244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e4e6f6465526566244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4d75742443244b24432456244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e496e7465726e616c24475424244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e45646765244754243130696e736572745f6669743137683061363937626335666465326231336145005f5a4e35616c6c6f633131636f6c6c656374696f6e733562747265653673656172636839315f244c5424696d706c2475323024616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e4e6f6465526566244c5424426f72726f77547970652443244b24432456244324547970652447542424475424313466696e645f6b65795f696e6465783137686536623733386637393339303364333045005f5a4e35616c6c6f633131636f6c6c656374696f6e733562747265653672656d6f76653235395f244c5424696d706c2475323024616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e48616e646c65244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e4e6f6465526566244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4d75742443244b24432456244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4c65616624475424244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4b562447542424475424313472656d6f76655f6c6561665f6b763137686636353666646236383034393666356645005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b244324562447542432356d657267655f747261636b696e675f6368696c645f656467653137683533393536653662353261323335336645005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b2443245624475424313662756c6b5f737465616c5f72696768743137683438363763626336383436386438373545005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b2443245624475424313562756c6b5f737465616c5f6c6566743137686265373332623332326366316630363345005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b244324562447542438646f5f6d657267653137686361323339646239313961656466353545002e4c706372656c5f6869323437002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e3731002e4c706372656c5f6869323438002e4c706372656c5f6869323530002e4c706372656c5f6869323439002e4c706372656c5f6869323531002e4c706372656c5f6869323533002e4c706372656c5f6869323532002e4c706372656c5f6869323534002e4c706372656c5f6869323535002e4c706372656c5f6869323537002e4c706372656c5f6869323536002e4c706372656c5f6869323538002e4c706372656c5f6869323539005f5a4e35616c6c6f6335626f7865643136426f78244c542454244324412447542431336e65775f756e696e69745f696e3137686638333630623536383435663835656545005f5a4e35616c6c6f6335626f7865643136426f78244c542454244324412447542431336e65775f756e696e69745f696e3137683561653632666364393337396638343545005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f646532313448616e646c65244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e4e6f6465526566244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4d75742443244b24432456244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e496e7465726e616c24475424244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e45646765244754243130696e736572745f6669743137686534333465396138336332386637346245005f5a4e35616c6c6f633131636f6c6c656374696f6e733562747265653673656172636839315f244c5424696d706c2475323024616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e4e6f6465526566244c5424426f72726f77547970652443244b24432456244324547970652447542424475424313466696e645f6b65795f696e6465783137683363626534356664313135636632613845005f5a4e35616c6c6f633131636f6c6c656374696f6e733562747265653672656d6f76653235395f244c5424696d706c2475323024616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e48616e646c65244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e4e6f6465526566244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4d75742443244b24432456244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4c65616624475424244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4b562447542424475424313472656d6f76655f6c6561665f6b763137686163343833363639623134363965653145005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f64653132354e6f6465526566244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4d75742443244b24432456244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4c6561664f72496e7465726e616c24475424313663686f6f73655f706172656e745f6b763137683737353737376565343533343639326445005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b244324562447542432356d657267655f747261636b696e675f6368696c645f656467653137683463636466393462393066383632383945005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b2443245624475424313662756c6b5f737465616c5f72696768743137683564316334326335313466346564393245005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b2443245624475424313562756c6b5f737465616c5f6c6566743137686632656564333962323432376663326445005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b244324562447542438646f5f6d657267653137683163656239623437396339613039313345002e4c706372656c5f6869323630002e4c706372656c5f6869323631002e4c706372656c5f6869323633002e4c706372656c5f6869323632002e4c706372656c5f6869323634002e4c706372656c5f6869323636002e4c706372656c5f6869323635002e4c706372656c5f6869323637002e4c706372656c5f6869323638002e4c706372656c5f6869323730002e4c706372656c5f6869323639002e4c706372656c5f6869323731002e4c706372656c5f6869323732005f5a4e34636f726535736c69636534736f727437726563757273653137683135373632303634376162396230656445005f5a4e34636f726535736c69636534736f72743235696e73657274696f6e5f736f72745f73686966745f6c6566743137686335633630633064646564353663303445005f5a4e34636f726535736c69636534736f72743134627265616b5f7061747465726e733137683666373839623434376138303465306245005f5a4e34636f726535736c69636534736f727432327061727469616c5f696e73657274696f6e5f736f72743137683166666132343636346439353362366245005f5a4e34636f726535736c69636534736f72743868656170736f72743137686335333661303961646638383239306245002e4c4350493136315f30005f5a4e35616c6c6f63377261775f7665633139526177566563244c54245424432441244754243136726573657276655f666f725f707573683137683432383261643562666265636465353945002e4c706372656c5f6869323733005f5a4e31387370617273655f6d65726b6c655f74726565356d65726765356d657267653137683435343932333464653765393762396445002e4c706372656c5f6869323736005f5a4e347574696c33736d7431316e65775f626c616b6532623137683834643333396363633032326665326245005f5a4e31387370617273655f6d65726b6c655f74726565356d6572676531304d6572676556616c756534686173683137683533636430316136373535316464336445002e4c706372656c5f6869323734002e4c706372656c5f6869323735005f5a4e31387370617273655f6d65726b6c655f74726565356d6572676531356d657267655f776974685f7a65726f3137683538623264626366313530366365656145002e4c706372656c5f6869323737002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e3331002e4c4350493136375f30002e4c4350493136375f31002e4c4350493136375f32002e4c4350493136375f33002e4c706372656c5f6869323738002e4c706372656c5f6869323739002e4c706372656c5f6869323830002e4c706372656c5f6869323831002e4c706372656c5f6869323832005f5a4e34636f726535736c69636534736f72743236696e73657274696f6e5f736f72745f73686966745f72696768743137686462656630303031353630316236376245002e4c706372656c5f6869323833002e4c4350493137315f30005f5a4e35616c6c6f63377261775f7665633139526177566563244c54245424432441244754243136726573657276655f666f725f707573683137683234396264636565353330343130653645002e4c706372656c5f6869323834005f5a4e39385f244c5424636b625f7374642e2e686967685f6c6576656c2e2e517565727949746572244c54244624475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137686531373133353834643233626333376245002e4c706372656c5f6869323835005f5a4e34636f726533707472373964726f705f696e5f706c616365244c5424636b625f7374616e64616c6f6e655f74797065732e2e67656e6572617465642e2e626c6f636b636861696e2e2e5363726970744275696c646572244754243137683631303764363938626431323933343345002e4c706372656c5f6869323838002e4c706372656c5f6869323836002e4c706372656c5f6869323837002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e3439002e4c706372656c5f6869323930002e4c706372656c5f6869323839002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e313133002e4c706372656c5f6869323931002e4c706372656c5f6869323932002e4c706372656c5f6869323936002e4c706372656c5f6869323933002e4c706372656c5f6869323934002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e3437002e4c706372656c5f6869323935002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e313138002e4c706372656c5f6869333030002e4c706372656c5f6869323937002e4c706372656c5f6869323938002e4c706372656c5f6869323939002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e313236002e4c706372656c5f6869333039002e4c706372656c5f6869333031002e4c706372656c5f6869333032002e4c706372656c5f6869333033002e4c706372656c5f6869333034002e4c706372656c5f6869333035002e4c706372656c5f6869333036002e4c706372656c5f6869333037002e4c706372656c5f6869333038002e4c706372656c5f6869333130002e4c706372656c5f6869333133002e4c706372656c5f6869333131002e4c706372656c5f6869333132002e4c706372656c5f6869333134002e4c706372656c5f6869333135002e4c706372656c5f6869333136002e4c706372656c5f6869333137002e4c706372656c5f6869333138002e4c706372656c5f6869333139002e4c706372656c5f6869333230002e4c706372656c5f6869333231002e4c706372656c5f6869333232002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3532002e4c706372656c5f6869333235002e4c706372656c5f6869333233002e4c706372656c5f6869333234002e4c706372656c5f6869333236002e4c706372656c5f6869333330002e4c706372656c5f6869333237007374722e32002e4c706372656c5f6869333238002e4c706372656c5f6869333239002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e3438002e4c706372656c5f6869333335002e4c706372656c5f6869333434002e4c706372656c5f6869333435002e4c706372656c5f6869333535002e4c4a54493138355f30002e4c42423138355f333137002e4c42423138355f323530002e4c42423138355f323537002e4c42423138355f323631002e4c42423138355f323733002e4c42423138355f323739002e4c706372656c5f6869333332002e4c706372656c5f6869333334002e4c706372656c5f6869333437002e4c706372656c5f6869333438002e4c706372656c5f6869333439002e4c706372656c5f6869333631002e4c706372656c5f6869333539002e4c706372656c5f6869333436002e4c706372656c5f6869333530002e4c706372656c5f6869333531002e4c706372656c5f6869333532002e4c706372656c5f6869333337002e4c706372656c5f6869333338002e4c706372656c5f6869333331002e4c706372656c5f6869333333002e4c706372656c5f6869333533002e4c706372656c5f6869333534002e4c706372656c5f6869333336002e4c706372656c5f6869333432002e4c706372656c5f6869333433002e4c706372656c5f6869333339002e4c706372656c5f6869333430002e4c706372656c5f6869333431002e4c706372656c5f6869333537002e4c706372656c5f6869333538002e4c706372656c5f6869333536002e4c706372656c5f6869333632002e4c706372656c5f6869333630005f5a4e397374616b655f736d7431315f42554444595f484541503137683461653061383139636232383364363745005f5a4e397374616b655f736d7431375f46495845445f424c4f434b5f484541503137683665376238383336646466636566323245002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3134002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3237002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3732002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3733002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3734002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3735002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3736002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3737002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3738002e4c6c696e655f7461626c655f737461727430002e4c6c696e655f7461626c655f737461727431006c69622e63002478002478002478002478002e4c32002e4c33002e4c3335002e4c3437002e4c3132002e4c3739002e4c3830002e4c3134002e4c3135002e4c3136002e4c3831002e4c3138002e4c3230002e4c3231002e4c3738002e4c3235002e4c3236002e4c3237002e4c3238002e4c3331002e4c3332002e4c3333002e4c3334002e4c3330002e4c3137002e4c3239002e4c3130002e4c313433002e4c313437002e4c313438002e4c313439002e4c323033002e4c313532002e4c323034002e4c313735002e4c313736002e4c313632002e4c323031002e4c313737002e4c313638002e4c313730002e4c313738002e4c313731002e4c313733002e4c313536002e4c313539002e4c313630002e4c313631002e4c313634002e4c323035002e4c313537002e4c313637002e4c313534005f5f636b625f7374645f6d61696e005f7374617274006d656d6d6f7665006d656d637079006d656d636d70006d656d73657400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000120000000000000060010100000000006001000000000000a00c00000000000000000000000000001000000000000000000000000000000009000000010000000200000000000000000e010000000000000e000000000000cc1600000000000000000000000000000800000000000000000000000000000013000000010000000600000000000000cc34010000000000cc240000000000005c5501000000000000000000000000000400000000000000000000000000000019000000010000000300000000000000289a020000000000287a010000000000a80000000000000000000000000000000800000000000000000000000000000020000000010000000300000000000000d09a020000000000d07a010000000000b80000000000000000000000000000000800000000000000000000000000000026000000080000000300000000000000889b020000000000887b01000000000000200800000000000000000000000000010000000000000000000000000000002b0000000100000000000000000000000000000000000000887b0100000000000c02000000000000000000000000000001000000000000000000000000000000390000000100000000000000000000000000000000000000947d01000000000078260000000000000000000000000000010000000000000000000000000000004500000001000000000000000000000000000000000000000ca401000000000020020000000000000000000000000000010000000000000000000000000000005400000001000000000000000000000000000000000000002ca601000000000050130000000000000000000000000000010000000000000000000000000000006200000001000000300000000000000000000000000000007cb9010000000000df4f0000000000000000000000000000010000000000000001000000000000006d00000001000000000000000000000000000000000000005b090200000000002c1c0000000000000000000000000000010000000000000000000000000000007d0000000100000000000000000000000000000000000000872502000000000024000000000000000000000000000000010000000000000000000000000000008d0000000300007000000000000000000000000000000000ab250200000000002b000000000000000000000000000000010000000000000000000000000000009f0000000100000000000000000000000000000000000000d625020000000000d71e000000000000000000000000000001000000000000000000000000000000ab0000000100000030000000000000000000000000000000ad440200000000002300000000000000000000000000000001000000000000000100000000000000b40000000200000000000000000000000000000000000000d044020000000000602301000000000013000000220c000008000000000000001800000000000000bc00000003000000000000000000000000000000000000003068030000000000ce00000000000000000000000000000001000000000000000000000000000000c60000000300000000000000000000000000000000000000fe68030000000000c466000000000000000000000000000001000000000000000000000000000000",
        "0x"
      ],
      "witnesses": [
        "0x550000001000000055000000550000004100000068d12bd305512c0feb84deaabd5ebddd6a514e1a7b54ac023e54064218ccbe156ad8ceac6e06465da09d3a925c6fe39c68a461a4b36fe51b74ea93e5db6680c800"
      ]
    },
    "0xbe3777fa551ec2de85ece9cca9918eefc953db190d52426d74c5f1cc73b2868c": {
      "version": "0x0",
      "cell_deps": [
        {
          "out_point": {
            "tx_hash": "0xf8de3bb47d055cdf460d93a2a6e1b05f7432f9777c8c474abf4eec1d4aee5d37",
            "index": "0x0"
          },
          "dep_type": "dep_group"
        }
      ],
      "header_deps": [],
      "inputs": [
        {
          "since": "0x0",
          "previous_output": {
            "tx_hash": "0xdfc4f59052fa596a2a8d0581be95450ce859e2da28c07aedb603d23429421f88",
            "index": "0x0"
          }
        }
      ],
      "outputs": [
        {
          "capacity": "0xec8d92f3e00",
          "lock": {
            "code_hash": "0x9bd7e06f3ecf4be0f2fcd2188b23f1b9fcc88e5d4b65a8637b17723bbda3cce8",
            "hash_type": "type",
            "args": "0x61a0d1fa2b4a4536a778659d5d87b88e82188b17"
          },
          "type": {
            "code_hash": "0x00000000000000000000000000000000000000000000000000545950455f4944",
            "hash_type": "type",
            "args": "0x89b5f5bcf25ed2a1b3486c8a2d6306f72ddd86c8788952dd17e1da1f8ea64a5b"
          }
        },
        {
          "capacity": "0xae968171180",
          "lock": {
            "code_hash": "0x9bd7e06f3ecf4be0f2fcd2188b23f1b9fcc88e5d4b65a8637b17723bbda3cce8",
            "hash_type": "type",
            "args": "0x61a0d1fa2b4a4536a778659d5d87b88e82188b17"
          },
          "type": null
        }
      ],
      "outputs_data": [
        "0x7f454c460201010000000000000000000200f30001000000e426010000000000400000000000000080750200000000000100000040003800050040001400120006000000040000004000000000000000400001000000000040000100000000001801000000000000180100000000000008000000000000000100000004000000000000000000000000000100000000000000010000000000e416000000000000e41600000000000000100000000000000100000005000000e416000000000000e426010000000000e426010000000000fa84000000000000fa8400000000000000100000000000000100000006000000e09b000000000000e0bb010000000000e0bb01000000000028010000000000002821080000000000001000000000000051e574640600000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007a740100000000008c740100000000009e74010000000000b674010000000000cc740100000000001695010000000000149501000000000018950100000000001c950100000000002095010000000000f674010000000000000000000000000001000000000000006486010000000000617474656d707420746f206164642077697468206f766572666c6f7700000000617474656d707420746f2073756274726163742077697468206f766572666c6f7700000000000000f67401000000000001000000000000000100000000000000308c01000000000008c9bcf367e6096a3ba7ca8485ae67bb2bf894fe72f36e3cf1361d5f3af54fa5d182e6ad7f520e511f6c3e2b8c68059b6bbd41fbabd9831f79217e1319cde05bf6740100000000000000000000000000010000000000000048800100000000000000000000000000617474656d707420746f207368696674206c6566742077697468206f766572666c6f7700000000000000000000000000617474656d707420746f206d756c7469706c792077697468206f766572666c6f77000000000000000000000000000000617474656d707420746f2073756274726163742077697468206f766572666c6f77000000000000000000000000000000617474656d707420746f2073686966742072696768742077697468206f766572666c6f77000000000000000000000000617474656d707420746f206164642077697468206f766572666c6f776c6561662073697a65206d75737420626520616c69676e20746f203136206279746573007c0301000000000023000000000000007265717569726573206d6f7265206d656d6f727920737061636520746f20696e697469616c697a65204275646479416c6c6f630000000000b00301000000000033000000000000006f7574206f66206d656d6f72790000000000000000000000617474656d707420746f20646976696465206279207a65726f00000000000000617474656d707420746f206164642077697468206f766572666c6f77427974655265616465724279746533325265616465724279746573526561646572000000617474656d707420746f2073756274726163742077697468206f766572666c6f775363726970745265616465725769746e65737341726773526561646572556e6b6e6f776e000000f67401000000000008000000000000000800000000000000a688010000000000456e636f64696e674f766572666c6f7776616c69646174654c656e6774684e6f74456e6f75676800f67401000000000008000000000000000800000000000000a6880100000000004974656d4d697373696e67496e6465784f75744f66426f756e6429426f72726f774572726f72426f72726f774d75744572726f7200000000b47701000000000018000000000000000800000000000000e680010000000000a28201000000000056830100000000002020202052656164446174612c0a2c20280a282c307830303031303230333034303530363037303830393130313131323133313431353136313731383139323032313232323332343235323632373238323933303331333233333334333533363337333833393430343134323433343434353436343734383439353035313532353335343535353635373538353936303631363236333634363536363637363836393730373137323733373437353736373737383739383038313832383338343835383638373838383939303931393239333934393539363937393839390000b477010000000000080000000000000008000000000000008e8301000000000098830100000000004e840100000000002829000000000000b477010000000000080000000000000008000000000000004e8601000000000054727946726f6d536c6963654572726f72636b622d64656661756c742d68617368616c726561647920626f72726f77656400000000000000f674010000000000000000000000000001000000000000004880010000000000616c7265616479206d757461626c7920626f72726f776564f67401000000000000000000000000000100000000000000368001000000000063616c6c656420604f7074696f6e3a3a756e77726170282960206f6e206120604e6f6e65602076616c75650000000000f67401000000000001000000000000000100000000000000308c010000000000617474656d707420746f206164642077697468206f766572666c6f77726561645f6174206069662073697a65203c20726561645f6c656e60726561645f6174206069662064732e63616368655f73697a65203e2064732e6d61785f63616368655f73697a6560726561645f617420606966206375722e6f6666736574203c2064732e73746172745f706f696e74207c7c202e2e2e60726561645f61742060696620726561645f706f696e74202b20726561645f6c656e203e2064732e63616368655f73697a656076616c69646174653a2073697a65203e206375722e736f757263652e746f74616c5f73697a65756e7061636b5f6e756d6265726765745f6974656d5f636f756e74636f6e766572745f746f5f753634636f6e766572745f746f5f7538636f6e7665727420746f205665633c75383e000000b691010000000000180000000000000008000000000000008a900100000000004669656c64436f756e744f75744f66426f756e64556e6b6e6f776e4974656d4f6666736574486561646572546f74616c53697a65436f6d6d6f6e0000000000000000000000000000617474656d707420746f206164642077697468206f766572666c6f770000000063616c6c65642060526573756c743a3a756e77726170282960206f6e20616e2060457272602076616c75650000000000f674010000000000100000000000000008000000000000006474010000000000f674010000000000000000000000000001000000000000006486010000000000617373657274696f6e206661696c65643a20636865636b706f696e745f646174612e69735f6e6f6e652829617373657274696f6e206661696c65643a207374616b655f61745f646174612e69735f6e6f6e6528290000000006000000000000000900000000000000060000000000000006000000000000000b000000000000000a000000000000000a000000000000000400000000000000080000000000000004000000000000002c0901000000000023090100000000001d0901000000000017090100000000000c090100000000000209010000000000f8080100000000009005010000000000e0040100000000008c050100000000001000000000000000017a5200017801011b0c02002c00000018000000161c0000181b000000440ed00d74810188028903920493059406950796089709980a990b9a0c9b0d1000000048000000fe3600000a000000000e0000100000005c000000f43600000a000000000e00001000000070000000ea3600000a000000000e00001000000084000000e036000008000000000000001000000098000000d436000008000000000000001c000000ac000000c83600004e00000000420e304a810188028903920493050018000000cc000000f63600003000000000420e20468101880289030010000000e80000000a370000080000000000000010000000fc000000fe36000008000000000000001000000010010000f236000008000000000000001000000024010000e636000008000000000000001000000038010000da3600000a000000000e0000140000004c010000d03600000e00000000420e10428101001800000064010000c63600005800000000420e4044810188020000001800000080010000023700005800000000420e404481018802000000180000009c0100003e3700005800000000420e40448101880200000018000000b80100007a3700005800000000420e40448101880200000014000000d4010000b63700005200000000420e404281010018000000ec010000f03700005800000000420e40448101880200000014000000080200002c3800005200000000420e40428101001800000020020000663800005800000000420e404481018802000000180000003c020000a23800004e00000000420e3044810188020000001c00000058020000d43800009a00000000420e2048810188028903920400000020000000780200004e390000dc00000000440e304c8101880289039204930594060000002c0000009c020000063a0000ee1a000000420ef0035a810188028903920493059406950796089709980a990b9a0c9b0d2c000000cc020000c45400001404000000420e80015a810188028903920493059406950796089709980a990b9a0c9b0d10000000fc020000a85800003c000000000e00001000000010030000d05800000a000000000e00001000000024030000c65800004c000000000e00001000000038030000fe5800004c000000000e0000100000004c03000036590000f4000000000e00002c00000060030000165a0000d403000000420eb00158810188028903920493059406950796089709980a990b9a0c00002c00000090030000ba5d0000f203000000420ec0015a810188028903920493059406950796089709980a990b9a0c9b0d20000000c00300007c610000d600000000420e504e81018802890392049305940695070018000000e40300002e6200004a00000000420e10448101880200000014000000000400005c6200003200000000420e10428101001800000018040000766200006e00000000420e5046810188028903001400000034040000c86200003400000000420e1042810100200000004c040000e46200006c00000000420e304c81018802890392049305940600000020000000700400002c6300006200000000420e304c81018802890392049305940600000010000000940400006a63000022000000000e000018000000a8040000786300003a00000000420e20468101880289030020000000c404000096630000fc00000000420e404e81018802890392049305940695070010000000e80400006e64000042000000000e000014000000fc0400009c6400009200000000420e104281010010000000140500001665000002000000000000001000000028050000046500003600000000000000180000003c050000266500007a00000000420e4044810188020000001800000058050000846500008200000000420e4044810188020000002400000074050000ea6500006001000000440ee00864810188028903920493059406950796089709100000009c0500002267000018000000000e000010000000b005000026670000040000000000000014000000c4050000166700000e00000000420e104281010010000000dc0500000c670000020000000000000014000000f0050000fa6600004201000000420e30428101002c0000000806000024680000e401000000420e705a810188028903920493059406950796089709980a990b9a0c9b0d001c00000038060000d86900005600000000420e304a810188028903920493050024000000580600000e6a00007803000000420e50528101880289039204930594069507960897090014000000800600005e6d00000e00000000420e10428101002400000098060000546d00007e01000000420e80015081018802890392049305940695079608000010000000c0060000aa6e0000120000000000000010000000d4060000a86e0000120000000000000014000000e8060000a66e00000e00000000420e104281010014000000000700009c6e00000e00000000420e10428101001400000018070000926e00007000000000420e90014281012c00000030070000ea6e0000bc01000000420e90015a810188028903920493059406950796089709980a990b9a0c9b0d140000006007000076700000b400000000420e10428101001400000078070000127100003800000000420e40428101001000000090070000327100000a0000000000000014000000a407000028710000b600000000420e104281010014000000bc070000c67100003a00000000420e404281010020000000d4070000e87100002001000000420ea0014e81018802890392049305940695071c000000f8070000e47200009800000000420e4048810188028903920400000014000000180800005c7300000e00000000420e10428101001000000030080000527300001600000000000000180000004408000054730000a200000000420e4046810188028903001400000060080000da7300007000000000420e90014281011c00000078080000327400005200000000420e304a81018802890392049305001800000098080000647400007c00000000420e5046810188028903001c000000b4080000c47400006200000000420e2048810188028903920400000010000000d408000006750000300000000000000018000000e8080000227500004c00000000420e1044810188020000001c00000004090000527500006800000000420e304a810188028903920493050018000000240900009a7500007c00000000420e5046810188028903001800000040090000fa7500005200000000420e204681018802890300180000005c090000307600005600000000420e10448101880200000020000000780900006a7600008201000000420e504e810188028903920493059406950700100000009c090000c8770000280000000000000010000000b0090000dc7700006200000000420e1018000000c40900002a7800006800000000420e30448101880200000018000000e0090000767800005400000000420e30448101880200000024000000fc090000ae7800007c01000000420e80015281018802890392049305940695079608970918000000240a0000027a00007800000000420e40468101880289030018000000400a00005e7a00007e00000000420e4046810188028903001c0000005c0a0000c07a0000a200000000420e50488101880289039204000000180000007c0a0000427b00007a00000000420e20468101880289030020000000980a0000a07b0000b200000000420e504c81018802890392049305940600000010000000bc0a00002e7c000010000000000000001c000000d00a00002a7c00007200000000420e5048810188028903920400000024000000f00a00007c7c0000ca02000000420ea0015081018802890392049305940695079608000010000000180b00001e7f000028000000000e0000240000002c0b0000327f00006401000000420ea0015081018802890392049305940695079608000024000000540b00006e8000007e05000000440e800864810188028903920493059406950796089709280000007c0b0000c48500001803000000420eb00256810188028903920493059406950796089709980a990b18000000a80b0000b08800009200000000420eb001468101880289032c000000c40b000026890000a003000000420ed0025a810188028903920493059406950796089709980a990b9a0c9b0d24000000f40b0000968c00008601000000420e90014c8101880289039204930594060000000000000000000002452c00014697000000e78000019308d00573000000130101932334116c2330816c233c916a2338216b2334316b2330416b233c5169233861692334716923308169233c91672338a1672334b167179600001306665c0ce208e6080c1306004013040040814597800000e78020d92338816205659b08458093050163080c09440146814601478147014873000000aa84630285080545638da406114463900418033b01631305004063786507854505445a8597600000e7800014aa8cae8a0c0c1306004097800000e78020e093020bc013850c402338516285659b88458093050163130600400943814601478147014873000000630d6510aa846309851011446397041083340163094463e29210a1a0014429a2054419a25a85814597600000e780600daa8cae8a0c0c5a8697800000e780a0d9114463708b023145b14b814597600000e780200b2a892e8a17e5ffff930515c691a003c51c0083c50c0003c62c0083c63c0022054d8d4206e206558e3364a600631a8b02214463788b0e3145b14b814597600000e780e0062a892e8a17e5ffff9305d5c131464a8597800000e780a0d285442da03145b14b814597600000e78040042a892e8a17e5ffff930535bf31464a8597800000e78000d08144da8923289120232a8121233c8120233031232334212323384123233c7123080c97500000e78040c20d4463870a00668597200000e780209eda8409a8014463870a00668597200000e780e09c2285a68597700000e780e0bf2a841315840361958330816c0334016c8334816b0339016b8339816a033a016a833a8169033b0169833b8168033c0168833c8167033d0167833d81661301016d828003c55c0083c54c0003c66c0083c67c0022054d8d4206e206558e3364a6001335840093753400b335b0004d8d15c531453149814597600000e78040f52a84ae8917e5ffff930535b03146228597800000e78000c18d4409bf63708b023145b14b814597600000e78060f22a892e8a17e5ffff930555ad65bd93592400fd190d4563f8a9023145b14b814597600000e780e0ef2a892e8a17e5ffff9305d5aa31464a8597800000e780a0bb91440d446dbd639ea908114691446685da85a28697500000e780e08b13f63500f199b306b5002338a120233cb1202330d1222334c12223389122130501630c0c97400000e780005d13050163da8597500000e780608a033901638334016423382121233c912009452330a122080c97500000e780c09b21cd31453149814597600000e78000e62a84ae8917e5ffff9305f5a03146228597800000e780c0b18d4459aa3145b14b814597600000e78060e32a892e8a17e5ffff9305559e31464a8597800000e78020af0d449144cdbb6380047605456380a47603360900833689006685da8597400000e780e07e13040002639e850e09456382a47403368900833609016685da8597400000e780c07c0544639e850e0d456385a47203360901833689016685da8597400000e780c07a2a86ae86080cb285368697400000e780607f8324012115456393a4100335816311c54a8597100000e780c0772d45636465016f10e00d93054bff0d456364b5006f10c00403c5dc0083c5cc0003c6ec0083c6fc0022054d8d4206e206558e83c51c0083c60c0003c72c0083873c00a205d58d4207e2075d8fd98d1147b366a600638ce50a03c55c0083c54c0003c66c0003877c0022054d8d42066207598e518d8d4563f6a56a7199c1456317b508080ce6855a8697400000e780e0684da8ae893145b14b814597600000e780a0ce2a892e8a17e5ffff9305e585314605a0ae892945a94b814597600000e780a0cc2a892e8a17e5ffff9305458329464a8597800000e7806098814403358163e30205c80335016397100000e780c06895b9032c4121033481218339012203398122033a0123833b8123c9bf93050bff0d45e377b57403c51c0183c50c0103c62c0103c73c0122054d8d42066207598e3367a600080ce6855a8697400000e78000570334012103360122281a9146a28597400000e780605c0335812111c5228597100000e78040617279b6642685814597600000e78040c12a84ae89ca85268697800000e780808d23388120233c312123309122130501630c0c97600000e780804103390163033481631305016313070002ca852286814697600000e780800103350163e30405720335016483358163033601632330a122233cb1202338c120880a0c0c97600000e780202b13050163930600025147ca85228697600000e78060fd03350163e30c056e0335016483358163033601632330a122233cb1202338c120a8120c0c97600000e7800027080c1306004013040040814597700000e78000752338816205659b08a581054562151307150093050163080c01468146814701487300000021c54944567511c5367597100000e7804050766511c5566597100000e780604f4a8597600000e780e0c7166511c5727597100000e780e04de38f0ab0668597100000e780004d01be033a0163130510406367aa0685450544528597600000e78040acaa892efa0c0c1306004097700000e780607893040ac0138509402338916285659b88a581131784030507930501631306004081468147014873000000833501633335a000b3b5b4004d8d21c9527529d94e8597100000e780a04599b75285814597600000e780c0a5aa892efa0c0c528697700000e7800072114463708a024545454c814597600000e78080a32a8bae8b17d5ffff9305355f91a003c5190083c5090003c6290083c6390022054d8d4206e206558e3364a600631a8a02214463788a084545454c814597600000e780409f2a8bae8b17d5ffff9305f55a45465a8597700000e780006b054d2da04545454c814597600000e780a09c2a8bae8b17d5ffff9305555845465a8597700000e7806068014d2328a121232ab121233c8120233041232334612323387123233c8123080c97400000e780c05a49445275e30205e64e8597100000e780803699bd03c5590083c5490003c6690083c6790022054d8d4206e206558e3364a6001335840093753400b335b0004d8d15c54545454b814597600000e780a0932a842e8a17d5ffff9305554f4546228597700000e780605f0d4d85bf63708a024545454c814597600000e780c0902a8bae8b17d5ffff9305754c21bf93542400fd140d4563f8a4024545454c814597600000e780408e2a8bae8b17d5ffff9305f54945465a8597700000e780005a114d0d44e1a0639ea408114691444e85d285a28697400000e780402a13f63500f199b306b5002338a120233cb1202330d1222334c12223389122130501630c0c97400000e78060fb13050163d28597400000e780c028033b01630334016423386121233c812009452330a122080c97400000e780203a29cd4545454b814597600000e78060842a842e8a17d5ffff930515404546228597700000e78020500d4d75a24545454c814597600000e780c0812a8bae8b17d5ffff9305753d45465a8597700000e780804d0d44114d268ab9b56302041405456302a41403360b0083368b004e85d28597400000e780201d99cd2a86ae86080cb285368697400000e780a021032d012115456316ad1209456309a41003368b0083360b014e85d28597400000e780a01999cd2a86ae86080cb285368697400000e780201e032d01211545631aad0e0d456300a40e03360b0183368b014e85d28597400000e780201699cd2a86ae86080cb285368697400000e780a01a032d01211545631ead0a0335816311c55a8597100000e780001393058aff0d45e377b52093054affe373b52003c5990083c5890003c6a90083c6b90022054d8d4206e206558eb366a60003c5d90083c5c90003c6e90003c7f90022054d8d42066207598e3367a600080cce85528697400000e780a000033501222aee49c503340121f2642685814597500000e780a06c2a8a2eeaa285268697700000e780e038a5a00145814509a80545854531a00945894519a00d458d4597500000e78040400000832d412103348121033a0122033b8122833b0123033c812303358163e30605cc0335016397100000e780c00575b917d5ffff1305c51f9305100297500000e780a0c20000014a0335812119c50335012197100000e780000363080a3a0d45f265e37cb55a03451a0083450a0003462a0083063a0022054d8d4206e206558e518d854529446318b554167593050002e31fb568d667014b02f603c5970183c5870103c6a70183c6b70122054d8d4206e206558e518d83c5d70103c6c70183c6e70103c7f701a205d18dc2066207d98ed58d82154d8daae303c5170183c5070103c6270183c6370122054d8d4206e206558e518d83c5570103c6470183c6670103c77701a205d18dc2066207d98ed58d82154d8d2aff03c5970083c5870003c6a70083c6b70022054d8d4206e206558e518d83c5d70003c6c70083c6e70003c7f700a205d18dc2066207d98ed58d82154d8d2afb03c5170083c5070003c6270083c6370022054d8d4206e206558e518d83c5570003c6470083c667003ee603c77700a205d18dc2066207d98ed58d82154d8d2af70d45aaff23300120130d1121930d9165080cac1b97600000e780a0dd034501218945630cb5246303051003459d0183458d010346ad018346bd0122054d8d4206e206558e518d8345dd010346cd018346ed010347fd01a205d18dc2066207d98ed58d82154d8d2334a16403451d0183450d0103462d0183463d0122054d8d4206e206558e518d83455d0103464d0183466d0103477d01a205d18dc2066207d98ed58d82154d8d2330a16403459d0083458d000346ad008346bd0022054d8d4206e206558e518d8345dd000346cd008346ed000347fd00a205d18dc2066207d98ed58d82154d8d233ca16203451d0083450d0003462d0083463d0022054d8d4206e206558e518d83455d0003464d0083466d0003477d00a205d18dc2066207d98ed58d82154d8d2338a16209a82334016423300164233c016223380162130501632c131306000297700000e780404b012519c1b27419aa130501630d46da8597400000e780400f03340163e301042e033581632af2833401642685814597500000e7802038aa8b2e8ca285268697700000e780600423387163233c816323309164130501659305016397600000e78040b80385ed008385dd0003c6cd0083340165230fa162a205d18d231eb16203c59d0083c58d0003c6ad008386bd0022054d8d4206e206558e518d232ca16203c51d0083c50d0003c62d0083c63d0022054d8d4206e20683c55d00558e518d03c64d00a20583c66d0003c77d00d18d834b8165c2066207d98ed58d82154d8d2338a162327511c5327597500000e780a0440305e1638315c16303268163833601632307a11e2316b11e2324c11eb6f3127511c5228597100000e780c0c87d556300ab56050b26f671bb294419b232756301051c0305e11e8315c11e0326811e9e76230ba11c231ab11c2328c11cb6e713051162ac033d4697700000e780e0f23275233ca16023007163080c930581610d4697500000e780006e033b0121e3010b2e0305712283056122034651222303a11aa205d18d2312b11a0345212283451122034631228306412222054d8d4206e206558e518d2320a11a0345a121834591210346b1218346c12122054d8d4206e2068345e121558e518d0346d121a2058346f12103470122d18d03048121c2066207d98ed58d82154d8d2aef327597500000e7806033130591182c0b3d4697700000e78080e75ae323048118130501630c030d4697500000e780e06203350163e30505240335016483358163033601632330a122233cb1202338c12028130c0c97600000e7804087130501630c03114697500000e780205f03350163e30005220335016483358163033601632330a122233cb1202338c120130501630c0c97600000e7806083ba7d7a768334016303370164080cee85a68697600000e78020ec0c0c13060002326597700000e780601f833581632a8491c5268597100000e78080ad5a7511c56e8597100000e780a0ac0dc45a8597500000e78000251304300319a01304b0065265630d05f2528597100000e78040aa6ff0cff2080c9146d285726697400000e78020a3833b0121833401222685814597500000e780c0082a842e8bde85268697700000e78000d5e38004168344040063070b00228597100000e78060a50335812119c50335012197100000e78040a4526511c5528597100000e78060a30545638aa4024944639b042e080c0546814597400000e78040c80345012163090510033581218335012297600000e78000c42a84e9a4130501650c0397100000e780a0b228130c0397100000e780e0a6130501630c0397100000e78080ab3a747a768334016303370164080ca285a68697600000e78060d813050002814597500000e78000fcaa8b2e8b0c0c1306000297700000e78020c80335816311c5268597100000e780e0985a7511c5228597100000e780009893050002054685445e8597700000e780e09f1375f50f13043004631e95029305000209465e8597700000e780209e1375f50f13044004631095028334016583350166268597600000e78080b92a841375f50f630c052063070b005e8597100000e780c091033581656300051e0335016597100000e7808090c1aa0305712183056121034651212307a11aa205d18d2316b11a0345212183451121034631218306412122054d8d4206e206558e518d2324a11a033581228305012303348121833401222338a162230cb1621305f11b93050163254697700000e78080b813558403230ba11a13550403a30aa11a13558402230aa11a13550402a309a11a135584012309a11a13550401a308a11a135584002308a11aa307811a13d58403230fa11a13d50403a30ea11a13d58402230ea11a13d50402a30da11a13d58401230da11a13d50401a30ca11a13d58400230ca11aa30b911a130501650c0397100000e780a0aa080c0c0397100000e78020840334016503360166833401210337012213050163a285a68697600000e780a0bb0335812111c5268597000000e780207e0335816511c5228597000000e780207d13050002814597500000e78040ddaa8d2e8b930501631306000297700000e78040a9a8030c0397100000e780c08d3e65fe6597600000e780c09f2a841375f50f05ed080cac03054697600000e780003e0345012105e10334812283340122080cac03094697600000e780403c0345012163020510034411215e6511c53e6597000000e780c07463070b006e8597000000e780e0731375f40f29c11a6597500000e78000ec6ff06fbb17d5ffff1305c5d9f1456ff02fed11456ff08fe863070b005e8597000000e78080700335816511c5268597000000e780806f1a6597500000e78000e8527511c54e8597000000e780006e567511c5367597000000e780206d766511c5566597000000e780406c4a8597500000e780c0e4166511c5727597000000e780c06a63870a00668597000000e780e06901446fe0dfcd3145da856ff02fe017d5ffff130525d297c5ffff9386255d09a817d5ffff130505d197c5ffff9386055c9305b002100c97400000e780403f00000335012283358122258da18d4d8d3d44e31a05ee080c2c13054697600000e780c032833b012263880b0c033581212af60335812283350123033681238336012136f22338a164233cb1642330c166aefbaaf7def3080c2c13094697600000e780c02e033c0122630b0c08033581212aee0335812283350123033681238336012136ea2338a164233cb1642330c1662334b1202330a120e2ff881397000000e780c0749374f50fa81b97000000e780e0731375f50f51446399a43c130501658c1397100000e7802082080cac1b97100000e780608103360166033501226313a602833501210335016597700000e780a0c7133a150001a80344012129b50344012149ae014a0335812119c50335012197000000e78080540335816519c50335016597000000e780605363000a36130581618c1397100000e7808080080c9305816197000000e780806f8335012241456397a54403350121834585002ee583459500aefc8345a500aef88345b500aef48345c500aef08345d5002efc8345e5002ef88345f5002ef4834505002ee183451500aeec83452500aee883453500aee483454500aee0834555002ef0834565002eec833581210346750032e889c597000000e780a0491305816197000000e780e0612ae613050165ac1b97000000e7802076080c9305016597000000e78020658335012241456394a53a03350121834585002ee2834495008345a500aef98345b500aef58345c500aef18345d5002ef98345e5002ef58345f5002ef183450500aefd83451500aeed83452500aee983453500aee583454500aee1834555002eed834565002ee983358121034a750089c597000000e780803f1305016597000000e780c0572afd1305016597000000e78080612a8d080c13060002ee8597600000e78020d10345012101c503441121d1aa8335812113852500636eb52a130460036311ad1c4a752205aa75c2050a7662066a682208ca68c208620a939284004e7342032e7462048e76b363d500d18d6e6e220ece66c2062e6762070e65b367a800b3641a01126533e5a20033646400b3e575006e763366ce00d98ec58f418d8215558e8217b3e8a50033e8c7000346811085428347810b6315560a62762206c276c206a274e2048273a20362634203c26ee20e667f220f467e420e267a620a0675b36fa600c58ee660a200466d420da665e205066533e7a30033e66e002a653364af003365ca01b3e6f6018a64b3e49000b3e5a501598e418d8216c58d0216c98e4d8e639857043337c800ba876384d800b3b7d8006395071c3275f265638aa50e3275f265c5a817d5ffff1305c59397d5ffff938645969305b002130601652db1639457083275f2656380a5023275f26531a83275f2656383a5043275f26589a01145f2656ff0af9d1275d26533b6a500631d0616127652673335c700b275f266b385b640898d3305c740b3c5b8003345a8004d8d1304700329e56da01275d2653337b500631907141277d26433359700b275f2679d8d898d33059740b58d318d4d8d1304a00311ed32756386a80032753335150121a01275333505011304800335c10335016597500000e78040970335816197500000e7808096628597500000e780e0955e8597500000e7804095a5b41275d265b3b7a500ede73385d840198db305c84012775266b334e600b276f267b386d740858e198e358db18d4d8d1304900345f10335016597500000e78020910335816197500000e7806090628597500000e780c08f5e8597500000e780208f014411b417c5ffff1305e57e97c5ffff93866503f9bc17c5ffff1305c57d97c5ffff9386c5089305b00213060163e9b417c5ffff1305257c97c5ffff938625074dbc17c5ffff1305057b97c5ffff9386050645b417c5ffff1305e5589305b0026ff02f8b17c5ffff1305e5ffc9ba17c5ffff130545016ff08f8917c5ffff130585006ff0cf8817c5ffff1305c5ff6ff00f8817c5ffff130505ff6ff04f8741456ff0ef8297300000e7808057000097300000e780a058000097000000e78060ff00001723000067002361173300006700e39d797106f422f026ec4ae84ee43284ae892a89328597200000e780e05eaa8405c163e38900a2892685ca854e8697600000e780e0334a8597300000e780009a2685a2700274e2644269a26945618280011106ec22e826e42a8497200000e780a05aaa8401c926858145228697600000e78020232685e2604264a2640561828017030000670023f717030000670023f717030000670023f717030000670083fb97000000e78080f40000411106e497300000e780a04b0000397106fc22f82a840a85194697500000e78040a702650dc14265a26502662af42ef032ec2c08228597500000e780a0cce27042742161828017c5ffff1305256397c5ffff938625ee9305b002300897400000e78060d10000397106fc22f82a840a851d4697500000e780c0a102650dc14265a26502662af42ef032ec2c08228597500000e78020c7e27042742161828017c5ffff1305a55d97c5ffff9386a5e89305b002300897400000e780e0cb0000397106fc22f82a840a85214697500000e780409c02650dc14265a26502662af42ef032ec2c08228597500000e780a0c1e27042742161828017c5ffff1305255897c5ffff938625e39305b002300897400000e78060c60000397106fc22f82a840a85354697500000e780c09602650dc14265a26502662af42ef032ec2c08228597500000e78020bce27042742161828017c5ffff1305a55297c5ffff9386a5dd9305b002300897400000e780e0c00000397106fcaa852800014697500000e7806091226519cd6265c26522662af82ef432f0081097500000e78000afe2702161828017c5ffff1305854d97c5ffff938685d89305b002101097400000e780c0bb0000397106fc22f82a840a85054697500000e780208c02650dc14265a26502662af42ef032ec2c08228597500000e78080b1e27042742161828017c5ffff1305054897c5ffff938605d39305b002300897400000e78040b60000397106fcaa852800094697500000e780c086226519cd6265c26522662af82ef432f0081097500000e780e09ce2702161828017c5ffff1305e54297c5ffff9386e5cd9305b002101097400000e78020b10000397106fc22f82a840a85154697500000e780808102650dc14265a26502662af42ef032ec2c08228597500000e780e0a6e27042742161828017c5ffff1305653d97c5ffff938665c89305b002300897400000e780a0ab0000797106f422f02a840a85194697400000e780007c026519c94265a265026608e80ce410e0a27002744561828017c5ffff1305a53897c5ffff9386a5c39305b0021306f10197400000e780c0a60000011106ec22e826e44ae02e892a84130505041306800b814597600000e780c0ec17c5ffff930505c213060004228597600000e78040f813053900a14522868346e5ff0347d5ff8347f5ff83440500a206d98ec207e204c58f0347150083442500dd8e834735000217a214458fc217830445005d8f1c62d98ee214c58ebd8e14e2fd1521062105c5fd0345090068f4e2604264a26402690561828069ce797106f422f026ec4ae84ee452e03284ae842a89687193050008b389a54063f6c9082330090e130a09065295a6854e8697600000e78040330335090493050508033689042330b904133505f81345150032952334a9044a85d28597000000e78000083304344113051008ce94636fa402930900080335090493050508033689042330b904133505f81345150032952334a9044a85a68597000000e7804004130404f893840408e3e789fc0335090e4a9513050506a685228697600000e780c02a0335090e22952330a90ea2700274e2644269a269026a45618280417186f7a2f3a6efcaebcee7d2e356ff5afb5ef762f366ef6aeb6ee72e892a842801130600082401814597600000e78040d40d0941458345e9ff0346d9ff8346f9ff03470900a205d18dc206620703461900d98e03472900d58d0216834639002217598e03074900c216558ed18d6217d98d8ce07d15a104210955fd280213060004a28597600000e78080db2c603064833204053267b2772a65aae89776000083b4663d033884053e972a97a58db98d9774000083b4a43c93d605028215d58d338e9500b346fe004a652ae193d78601a216dd8e2a973303d700b345b30013d70501c215b3e8e500469eb345de0093d6f50386055267d274ea67bee41775000003356538b3ebd50026973e97318d398d9775000083b5a537135605020215518daa95ad8c8a7636f813d68401a214d18c3386e600330996003345a900935605014215b36cd500338abc0033459a009355f5030605f26672772a769774000083b48433b369b500ba96b296328c32f433c59200358d9774000083b464329357050202155d8daa94258fca752eec935787012217d98fae96b382f60033c5a200935605014215b36dd500ee94a58f13d5f703860792761666ea75aefc177700000337872e33eba700b296ae963345e800358d177700000337a72d9355050202154d8d2a97398e8e67bef0935586012216d18dbe96b383b60033c5a300135605014215518d2a97b98dae6a13d6f5038605d18d56934e933345a300135605020215498eb29433c53401ce69935685012215c98e338569004ee8b30ed50033c6ce00935706014216336df600b3009d0033c6d0006e6f9356f6030606b36fd6007a99fae033032b01b347130193d407028217c58f3e97b34467010e75aaf493d88401a21433e61401b3086500b298b3c7f80093d40701c21733e39700330be3003346cb002e75aaf81357f6030606b364e600aa92ae9233c69201135706020216598e329eb345be004e7913d78501a2154d8fb30559004af03388e5003346c800935206014216b36256003386c201318fee751355f7030607336ea700ae93ae86aeecde9333c5b301935d050202153365b501b30c4501b3cd7c01926793d58d01a21db3e5bd00be933e873efcb38db30033c5ad00935305014215336a750033059a01a98d93d7f5038605dd8db69eae9eb3c76e0093d607028217dd8e3696b18d93d78501a215dd8db387ee01b38eb700b3c6de0093d70601c216b3e3f6003383c300b345b30013d6f5038605b3ecc500e298fe98b3c5120113d605028215d18d2e953346f501935686012216d18e56e4338658013696b18d93d70501c215b3e8f500b382a80033c5d2009355f50306054d8d4e982698b3450a0193d605028215cd8eb690b3c5900093d78501a215cd8fb3050701b38ff500b3c6df0093d40601c21633e89600c290b3c6f00093d7f6038606d58fca9df29db3c6ad0193d406028216d58c338f6401b346cf0113d78601a216558fe676ee96338ae600b3449a0093d50401c214c58d2e9f3347ef009354f7030607d98c8a66b69eaa9eb3c5be0013d705028215d98d33871500398d935685012215c98e467b33856e01b30ed500b3c5be0013d50501c215b3eba500338deb00b346dd0013d5f6038606b3e0a600466c62963e96334576009355050202154d8d2a9fb345ff0093d68501a215d58d266e7296b309b60033c5a900935605014215558d2a9fb345bf0093d6f5038605b3edd5002676b29fa69fb3c51f0193d605028215cd8e3693b345930093d48501a215cd8c8675fe95b3839500b3c6d30093d70601c216d58f3e93b346930093d4f6038606b3e8960062673a9a669ab3460a0193d406028216c58eb692b3c4920193d58401a214c58d4279b3044901b38fb400b3c6df0093d40601c21633ea9600b3045a00a58d93d6f5038605d58db29eae9e33c5ae00935605020215c98eb382660033c5b200935585012215c98d33855e01b30cb500b3c6dc0013d50601c216b3eea600f69233c5b2009355f50306053363b50033063b010696b18f13d5070282175d8d3388a400b345180093d68501a215d58d62962e96318d935605014215b360d50006983345b8009355f50306054d8dba93ee93b3457a0093d605028215cd8eb387a601b3c5b70113d78501a215b3e4e500b385c301338a9500b346da0013d70601c216b3e3e6009e97bd8c93d6f4038604c58ee275ae9fc69fb3c47f0113d704028214458f3a9fb3441f0193d58401a214c58d827bde9fae9f33c7ef00935407014217458f3a9fb345bf0093d4f503860533ec95008665ae9caa9c33c7ec00935407020217458fba973d8d935485012215c98ce669338599012695298f935807014217336b1701b30cfb0033c79c009357f7030607b36df700ca8a4a96b305d60033c7be009357070202175d8fb307ef00bd8e93d48601a216c58e66762e96338dc6003346ed00135706014216b36ee600338efe00b346de0013d7f603860633efe6000676329a629a33471a00935407020217458fba92b3c5820193d48501a215cd8c8a68b3854801338a95003347ea00935707014217336cf700e292b3c7920093d4f7038607b3e097004267ba9f9a9fb3c77f0093d407028217c58f3e98b344680093d68401a214c58e2279ca9fb69fb3c7ff0093d50701c217dd8db3870501bd8e93d4f6038606c58e329536953346d501935406020216458e33085600b346d80093d48601a216c58e3a953695298e935406014216336396001a983346d8009356f6030606b362d600569d6e9d3346ac01935606020216d18eb69733c6b701135786012216598e3387a801b30ac700b3c6da0093d40601c216b3e39600b38df30033c6cd009356f6030606558e5e9a7a9ab3c5450193d605028215cd8eb3889601b3c5e80193d78501a215cd8fc675d295338ab700b346da0093d40601c21633ef9600fa98b3c7f80093d4f7038607c58fa675ae9f869fb3c66f0193d406028216d58cb38ec401b3c61e0093d58601a216d58db3863f01b38fb600b3c49f0093d60401c214c58eb69eb3c5be0093d4f5038605c58da66b5e953307c500b98e93d406028216c58eb69833c6c800935486012216458e66753a953295a98e93d40601c21633ec9600b30c1c0133c6cc009356f6030606336ed600e26833871a013e9733466700935606020216558e3303d601b346f30093d78601a216dd8e866a5697330dd7003346cd00135706014216598e3293b346d30013d7f6038606b3e0e600ca894a9a2e9ab3467a0013d706028216d98e3698b345b80013d78501a215d98dc66433079a00b38ee500b3c6de0093d70601c216dd8e3698b345b80093d7f5038605b3e3f5006279ca9f969fb3c5ef0193d705028215cd8fbe9db3c55d0013d78501a2154d8f226bb305fb01338fe500b347ff0093d50701c217dd8dae9d33c7ed009357f70306075d8fc2673e953a95298e9357060202165d8e32983347e8009357870122175d8f2695b307e5003d8e135506014216b362a60016983345e8001356f5030605518d2ae8469d729d33c5a601135605020215498eb29d33c5cd01935685012215c98e06756a95330dd5003346cd00135706014216b36fe600338ebf013346de009356f6030606d18ede9e869eb3c5d50113d605028215d18db388950133c61800135786012216598e33873e01b30dc700b3c5bd0093d40501c215b3ee9500f698b3c5c80013d6f50386054d8e569f1e9fb3458f0193d405028215cd8c2693b345730013d58501a2154d8db3052f01b383a500b3c4930093d50401c214c58db3846500258d1357f5030605498f6665aa97b697bd8d13d5050282154d8daa98b3c5d80093d68501a215d58d8a66be96b380b60033c5a000935705014215336af500b30b1a0133c5bb009355f50306053363b50026794a9d329d33c5a201935505020215c98db388b40033c5c800135685012215498e467c33058d01330fc500b345bf0093d70501c215cd8fbe98b3c5c80013d6f5038605b3e2c500667dea9dba9db3c5fd0113d605028215d18d2e983346e800135786012216518f33866d01da89b30ce600b3c5bc0093d40501c215c58d2e983347e8009354f7030607b36f9700c27dee934265aa9333c7d301935407020217d98cb38ac40133c7aa00135587012217598d027e33077e00b30ea700b3c49e0013d60401c214d18c33865401318d9356f5030605558da666b690aa90b3c6f00093d706028216dd8eb38a060133c5aa009357850122155d8db3878001aa97bd8e13d70601c21633e8e600c29a33c5aa009356f5030605b363d5006a9f1a9f33c5e501935505020215c98d2e9633456600935685012215c98e06657a95330dd500b345bd0013d70501c21533e3e500330fc300b345df0013d6f5038605d18d4665aa9c969c33c69401935606020216558eb29bb3c65b0013d78601a216558fb3862c013309d7003346c900935406014216336b9600da9b33c6eb001357f6030606598ece9efe9e33c74e01935407020217d98ca69833c7f801935687012217d98e3387be01330cd700b3449c0013d70401c214458fb3041701a58e13d5f6038606c98e2275aa97ae973d8f135507020217598db30f7501b3c5bf0013d78501a215d98df297338ab7003345aa00135705014215b362e500969f33c5bf008e689355f5030605b369b500469d329d33450d019355050202154d8db30e950033c6ce00ca7d135786012216598eb384ad01338dc4003345ad00135705014215498fba9e33c6ce00926c9357f6030606b36bf60066993699334669009357060202165d8eb29ab3c6da0093d78601a216dd8ee667ca97338ed7003346ce00135506014216518daa9a33c6da009356f60306063369d6008a652e9c1e9c33468b01935606020216d18e369f33467f004e68935786012216d18f33060c01338bc700b346db0013d60601c216558eb306e601b58fae7493d5f7038607dd8dd294ae94258f9357070202175d8f330f5701b3c5e50193d78501a215cd8fb385b401338cb70033478701935407014217336a9700529f33c7e701ca679354f703060733639700ea97ce973d8d135705020215598db303d500b3c6790013d78601a216558fb3869701b30cd70033459501935705014215b369f500ce93334577006e779357f50306055d8d72975e97398e9357060202165d8eb29fb3c7fb014e7e93d48701a217c58f7297338de7003346a601135706014216b36ae600d69f33c6f7012a779357f60306065d8e5a974a97b3c5e20093d705028215cd8fbe9eb345d901ee6693d48501a215cd8cb305d700b382b400b3c7570093d60701c217dd8eb69e33c7d401aa679354f7030607d98ce297aa97bd8e13d706028216d98eb69f3345f501135785012215598dc697330cf500b3c6860113d70601c21633e9e6004ae3ca9f3345f501ea761357f5030605b36be500e696b2963345da00135705020215598d330ad501334646018a7e135786012216598ef696b30dd6003345b501935605014215558d2a9a334646019356f6030606336bd600429d269d33c6a901935606020216558e329fb3c6e401ea6493d58601a216d58db3069d00b38cd50033469601935406014216458e329fb3c5e501ae6493d7f5038605b3e9f500a6929a92b3c55a0093d705028215cd8fbe93b34573008e7493d68501a215cd8eb3859200b38ab600b3c7570193d50701c217dd8db3877500bd8e13d7f6038606d98e629e369e3345c501135705020215598db302e501b3c6560013d78601a216d98e269e338cc60133458501135705014215b363e5009e9233c556009356f5030605336fd5007af6ee98de9833451601135605020215518d3303f50033c66b00ee76135786012216598ec696b30bd60033457501935605014215336ed5007293334566002e769356f5030605558d66965a96b18d93d605028215d58db386f5013347db00ca67935487012217d98c3e96338bc400b3c5650113d60501c215b3efc500fe96b58c93d5f4038604b3ecb400d69ece9eb345d90113d605028215d18d2e9a33c64901935486012216d18c33860e01b38ac400b3c5550113d60501c215d18d2e9a33c64401ca741357f6030606598ee294aa94a58d13d705028215d98dae96358d2a679357850122155d8d2697330de500b3c5a50113d70501c215b3eee50076e3b388de0033451501126c9356f50306053369d500e29be69b33c57301935605020215c98eb383460133c57c002a77935785012215c98f3385eb00338aa700b3c6460113d70601c216558fba93b3c677002e6893d7f6038606b3ebf600429b329bb3466e0193d706028216d58fbe9233465600ea75935686012216558eb306bb00330bd600b3c7670113d50701c2175d8daa92334656006a6e9357f6030606b369f600f29afa9a33c65f01935706020216d18f3e9333466f00ee66935486012216d18c3386da002696b18f93d60701c217dd8e3693b3c7640093d4f7038607c58fea95be952d8f935407020217d98ca69233c75700935787012217d98fe295b38ab700b3c4540193d50401c214b3efb400fe92b3c5570093d7f503ee74860533eff5007af6d294ca94258d935505020215c98d2e9333456900ce67135785012215498f3385f400330ca700b3c5850193d70501c21533eaf5005293b34567000e7793d7f5038605cd8f5a975e97b98e93d506028216d58dae98b3c61b018a7413d58601a216558d2697b304e500a58d93d60501c21533e9d500ca9833451501aa659356f5030605558db295ce9533c6be00935606020216558eb293b3c6790013d78601a216d98ec2953388b60033460601135706014216598eb293b3c676002e7793d5f6038606d58d56973e97398e935606020216558eb298b3c6170193d78601a216d58fb306c701b389d70033463601135706014216b36ee60076e3f69833c617014e779357f6030606336bf60062972a9733c6ef00935706020216d18fbe93334575008e6f135685012215518d3306f701330cc500b3c7870113d70701c2175d8fba93334575004a6e9357f5030605b36af500f294ae9433459a009357050202155d8daa92b3c555002a7a13d68501a215d18dd294b38c950033459501135605014215336dc500ea92b3c555006e6693d6f5038605b3ebd50032987a98b345090193d605028215cd8eb3846600b3459f004a7393d78501a215cd8fb30568003389b700b3c6260193d50601c216d58dae94a58f93d6f7038607dd8e4e963696318f9357070202175d8f33085700b3c60601ea6713d58601a216558d3e96b30dc5003347b701135607014217b369c7004e98334505011356f5032e670605336fc5007af662975a973345ed00135605020215518db302950033465b009357860122165d8e5297330be60033456501135705014215336ae500d292334556001356f5030605518de69fd69fb3c5f50113d605028215d18d3387150133c6ea00ea74935786012216d18f33869f00b38fc700b3c5f50193d40501c215b3e895004697b98f93d5f7038607dd8d4a9e5e9eb3c7ce0193d407028217c58fbe93b3c47b0013d68401a214458e7293b30e6600b3c7d70193d40701c217c58fbe933346760092649356f6030606558eee94aa94a58f93d607028217dd8e3383e600334565000e779357850122155d8d2697b30be500b3c6760193d70601c21633eef60072e3729333456500ce669357f50306053369f500da96ae9633c5d900935705020215c98fbe9333c57500ee75935485012215c98c3385b600338ba400b3c7670193d50701c217dd8dae93b3c674008a7a93d7f6038606b3e9f600d69fb29fb346fa0193d706028216dd8e369833460601ae77935486012216458efe97330cf600b3c6860193d40601c216c58e369833460601ce741355f6030606336aa600a69efa9e33c5d801135605020215518daa9233465f002a67935486012216458eba9e330fd6013345e5019357050142155d8daa92334656009357f60306065d8e5e973297b98d93d705028215dd8d2e9833460601ca67935486012216d18c3306f700b38cc400b3c5950113d70501c215b3efe5007e98b3c5040113d7f503ea678605b3eee50076f6da97ca97bd8e93d506028216cd8eb3885600b345190113d78501a2154d8fb3855701330bb700b3c6660193d70601c216b3eaf600d69833471701aa779354f7030607458fe297ce973d8d935405020215458d2a93b3c46900ca7693d58401a214c58dbe96b38bd500334575019356050142153369d5004a9333c56500ea759356f5030605c98efa95d2953345be00935405020215c98ca69333457a008e67135685012215498e3385f500330ca600b3c4840193d50401c214c58db38775003d8eae629354f6030606458e969cba9cb3c5950193d405028215c58db3836500334777004e63935487012217458fb3846c00330d9700b3c5a50113d50501c21533efa500fa9333457700ee6c9355f5030605b369b500669b369b33c56f019355050202154d8daa97bd8e8e7513d78601a216d98eda95338bb60033456501135705014215498f330ef70033c5c601ae769357f5030605336af500de96b29633c5da009357050202155d8d2a9833460601ce7f935786012216d18f3386f601b38bc70033457501935605014215558d2a98b3c50701ee7793d6f5038605b3ead5003e9c769cb345890193d605028215d58dae98b3c41e01926613d68401a214458eb304dc0033099600b3c5250193d40501c215c58dae98334616019354f6030606458eea97b2973d8f935407020217458f3a9833460601935486012216458ee697330cf60033478701935407014217b36e97007698334606011357f6030606aa74598e7ae332f6da94ce94258d135605020215518d3306150133c7c900935787012217d98f33875400b389e70033453501935405014215b36895004696b2ea3d8e1355f6030606b367a6005e93529333c565009355050202154d8daa93b3457a0013d68501a215d18d3306d3003383c50033456500935605014215b362d500969333c575009355f5030605b366b500ca9fd69f3345ff01935505020215c98d2e9e33c5ca01ea74135685012215498e33859f00330fa600b3c5e50193d40501c215cd8c269eb345c6014a6613d5f5038605c98d62963e96b18c13d504028214458daa93b3c77700ae7413d78701a2175d8f26963a9632e6318d135605014215518d2ae31e95aaee398d1356f5032a670605518d2afa4e97369733c5ee00135605020215518d2a9e33c6c601ea669357860122165d8eba96b29636ea358d935605014215558daaf67295aaf2318d1356f5038e760605518d2afe9a96ae9633c5d800135605020215518d2a98b3c505010e6613d78501a215d98d36962e9632ee318d135605014215518daafa4295aae62d8d9355f50306054d8daae23275ca75aa95fa9533c6b200d666135706020216598eb296358d0a779357850122155d8dba95aa952ef2b18d13d60501c215d18daefeb695aeea2d8d9355f5030605c98da8022ef6a1451060833605fc1861358e398e10e0fd1521052104f5f5be701e74fe645e69be691e6afa7a5a7bba7b1a7cfa6c5a6dba6d7d618280197186fca2f8a6f4caf0ceecd2e8d6e4dae05efc62f866f46af06eec906103bc8500329c636fcc34aa8988699376f50093b616003337a000f98e6380063a814a89466368d5008d462a87850a0581e3ede6fe83cb85013285d68597000000e780a03b6365ac322a8d1305000463f5aa323305ac4133555501814c89456368b5008d452a86850c0581e3edc5fe938d2c0063ea9d316145b3b5ad02639a0530b384ad02ea9463eaa43113893c006a847d19268a630d0902630c0d24233044015285639b0b00130600105285814597400000e780401b0860610408e1c10408e5e3f844fd17a5ffff13052502a5ac4ee0638b0d2e014b13098d0093891c005a85ee8597000000e780a03563030d201d05935435002330490163990b0052858145268697400000e7800016d29463e24425638669016109050b268ad1b7094963e72d0593098d02330a904105442285ee8597000000e780c0301d05135b350023b0990063990b00268581455a8697400000e780601133856401636195200504b3058a00e109aa84e39325fd11a02685d68597000000e7806028636fac2463860d262a8b938bfdff2a84638b0b161385edff9305f00363eda520854c5a846ae86ee463080d14aa843395ac00331d55013309a401636589186145b38da402c265ae9d3385ab022e9593098500130a0501636f2c0d03b50d000c612300b40013d68503a303c40013d605032303c40013d68502a302c40013d605022302c40013d68501a301c40013d605012301c400a181a300b40093558503a307b400935505032307b40093558502a306b400935505022306b40093558501a305b400935505012305b40093558500a304b4002304a4000c6180e500e15a85d6852686a28697000000e780c022058915ed5a85d6855e86a28697000000e780802183b5090013563500b295838605001d893395ac00c98e2380d50083350a00b29503860500518d2380a5004a846a99e37489f249a82685a26597000000e780c0185a85d6852686a28697000000e780801c83b58d0013563500b295038605001d893395ac00518d2380a50081cc1385f4ffa68b426de31c0dea97200000e780e0af0000426da26d63638c0a33058c40826523b0650123b4850188e923bca50123b0b50323b45503e6704674a6740679e669466aa66a066be27b427ca27c027de26d0961828017a5ffff1305a5daf14597200000e780a08e000017a5ffff130565d9f5b717a5ffff1305c5d8cdb717a5ffff130525d8e1bf17a5ffff130585d1ada817a5ffff1305e5d393054002c9b717a5ffff130505d65dbf17a5ffff130565cca1a817a5ffff1305c5d44db717a5ffff130525ce91a017a5ffff130585c79305300271b717a5ffff1305a5d629a85285d68597000000e780c002637bac0017a5ffff130585d997000000e7804005000017a5ffff1305e5c99305100289bf01cd1306000463f0c5027d153355b50005053315b500828017a5ffff130585c79305100239a017a5ffff1305a5c99305400297200000e7808080000097100000e780a00f000063efa5006382a5021345f5ffaa951305000463f2a50205453315b500828017a5ffff1305c5c229a017a5ffff130525c29305100239a017a5ffff130545bb9305300297100000e780207b000063e0a6041307f003636cc7001307000463fde500898e33d5c6003355b500828017a5ffff1305e5c029a017a5ffff130545c09305400297100000e7802077000017a5ffff130565cbb545f5b790659461137806fc3698636bd80c98699355660063e3e500ba8594e2094694e6b68763ebc508fd1593d8860393d2060313d3860293d3060213de860193de060113df8600b68736863e879387070463efe7062380c70013578603a383e700135706032383e70013578602a382e700135706022382e70013578601a381e700135706012381e7002182a380c7002384d700a387170123875700a386670023867700a385c7012385d701a384e70190621ce6fd159ce23e86c9f99385070463e7f50214e1233405010ce914ed828017a5ffff130565b4f14597100000e7806068000017a5ffff130525b3f5b717a5ffff130585b2cdb7717106f522f126ed4ae94ee552e1d6fcdaf8def4e2f0e6eceae82a841305000497550000138ae53e63718504175500009304253e8860631e05348864fd558ce063130512c870cc6cd068d464aae4aee032fc36f80a850c1897000000e780209c054588e413850401c5a803350a04631b053203358a04fd552330ba041ded03350a0883358a0703360a07aae02efc32f80a850c1897000000e78080e705452334aa040265a2654266e2662338aa04233cba042330ca062334da0603398a0663000902033509000c6110650ce20c6510610ce6130b0a04630825032a8991a403390a0603358a056373a902130509046368252983350a042330aa0685052330ba046315092209a823340a0619ac03350a0405052330aa0403350a00631e052803358a00fd552330ba001ded03350a0a83358a0903360a0983368a08aae4aee032fc36f80a850c1897000000e780408d05452334aa0013050a018a851306000397400000e780a0c083398a031305f003636335210545814c3315350163788500850c63840c1c0605e36c85fe83350a0363e3bc00e68503358a020146e146b386dc02aa96138406fdb385bc406389c516630d051c147803b9060061047d16e307d9fe033509008335890088e1033589008335090088e5047017550000130b852303350b0183358b03934af6ffe69a5686ca8697000000e78000cd93553500a695038605001d89854b3395ab00518d2380a50063f85c11130c000417550000130b651f138afaff63778a1333954b01b3143501ca9463e72413033d840203350b0183358b035686ca8697000000e780a0c793553500ea95038605001d893395ab00518d2380a500833a840003350b0183358b035286ca8697000000e780c0c493553500d695038605001d893395ab00518d2380a50008600c612380b40013d68503a383c40013d605032383c40013d68502a382c40013d605022382c40013d68501a381c40013d605012381c400a181a380b40093558503a387b400935505032387b40093558502a386b400935505022386b40093558501a385b400935505012385b40093558500a384b4002384a4000c6184e504e12114d28ae3e54cf119a00149528b03350b0005052330ab004a85aa700a74ea644a69aa690a6ae67a467ba67b067ce66c466d4d6182801795ffff1305657d21a81795ffff1305c5709305300231a01795ffff1305e57bf14597100000e780e02f00001795ffff1305a56ef9bf1795ffff1305057acdb797100000e780e049000017a5ffff1305d5b09795ffff9386c56915a017a5ffff1305b5af9795ffff9386a56809a817a5ffff130595ae9795ffff93868567c1450a8697100000e780e0440000317106fd22f926f54af14eed52e956e55ae1defce2f8e6f4eaf0eeec97550000938ce50183b50c04639d05382a8903b58c04fd5523b0bc041de9175500001304050048602c7c3078aae4aee032fc28002c1897000000e78060ae054528e42265c2656266827628e82cec30f034f403b50c0583b58c053335a9001345f5ffb335b9006d8d51c517550000130545fb2c75638e052090612300c90093568603a303d900935606032303d90093568602a302d900935606022302d90093568601a301d900935606012301d9002182a300c90013d68503a307c90013d605032307c90013d68502a306c90013d605022306c90013d68501a305c90013d605012305c90013d68500a304c9002304b900906165a203b50c0483b50c00050523b0ac04639b052a03b58c00fd5523b0bc0015ed175500001304c5f048704c6c50685464aae8aee4b2e036fc28002c1897f0ffffe780c04f054508e4130504012c001306000397400000e780408383ba0c03638f0a2283b98c02138afaff13848902854463809a04638b0922033b040003b50c0183b58c032686ca8697000000e780609593553500da9583c505001d8933d5a50005898504610469d5f91463e6440139a263030a108144930a0004268b63e49a00130b000483bb8c0303bc0c0161453385a4024e9513048502054d03b50c0183b58c032686ca8697000000e780808f638e091a833504fe13563500b2950386050093767500b316dd0093c6f6ff758e2380c500937515003306b040833604fe13661600329513563500369603460600937675003356d600058a51e2630b9b1263fe5b1333159500331575016295636e85131061146590e21065146190e691c12a89833d040003b50c0183b58c0385042686ca8697000000e780c08693553500ee95038605001d893315ad001345f5ff718d2380a5006104e3129af4d28405a023302901930585064a862334260123b02501930c050451a8638a090e814461453385a4024e9508610c612300b90013d68503a303c90013d605032303c90013d68502a302c90013d605022302c90013d68501a301c90013d605012301c900a181a300b90093558503a307b900935505032307b90093558502a306b900935505022306b90093558501a305b900935505012305b90093558500a304b9002304a9000c6123b425012330250103b50c00050523b0ac00ea704a74aa740a79ea694a6aaa6a0a6be67b467ca67c067de66d296182801795ffff1305c53029a01795ffff130525309305300231a01795ffff1305453bf14597100000e78040ef00001795ffff1305053493051002edb797100000e780a00900001795ffff130595709795ffff9386852909a81795ffff1305756f9795ffff93866528c145300097100000e780c00500005d7186e4a2e026fc4af84ef452f056ec83ba050263800a0a2e8a2a898065b35954034e8597000000e780200b83340a002ae02ee402e863e335078145636e54031396350032950d466370560983c6140003c70400a206d98e03c7240083c7340033045441d6944207e2075d8fd98e14e185052105e37a54fd2ee8226502662338b9002334a9002330c900a6600664e2744279a279027ae26a616182800a8581454e8697000000e780e007c2650265e37954f9d9b71795ffff13054535e54597100000e78040de00001145d68597100000e780c0560000411106e422e02a840dc51355c4030de993351500131534008e0511c597d0ffffe780401caa8599e597d0ffffe780801d0000a1452e85a285a26002644101828097d0ffffe780a01c0000411106e497000000e780e002fd55fe1585056315b500a2604101828011e597d0ffffe780201a000097d0ffffe780e01800005d7186e4a2e026fc2e966374b600014591a82a8408659314150063639600b284914563e39500914493d5c40393b51500139634008e0501c914600e0536f0a14636f42af811a002f42800141097100000e780e069a265426591e508e004e47d557e150505a6600664e27461618280411106e4054697000000e780c0f8fd55fe1585056315b500a2604101828011e597d0ffffe7800010000097d0ffffe780c00e0000797106f422f026ec4ae84ee452e06365d7046366e604aa89b304d7403389d5002685814597100000e780606b2a842e8aca85268697300000e780a03723b0890023b4490123b89900a2700274e2644269a269026a456182803685ba8519a03a85b28597100000e780203e0000797106f422f026ec4ae84ee452e06363d604aa89b304d6403389d5002685814597100000e780e0642a842e8aca85268697300000e780203123b0890023b4490123b89900a2700274e2644269a269026a456182803685b28597100000e7800038000063e8c60063e9d500b385c640329582803285b68511a0368597100000e780e0350000011106ec22e826e42a8410690865ae846319a6002285b28597000000e78040ec10680860931536002e9504e1050610e8e2604264a26405618280397106fc22f826f44af04eec52e856e4114a32892a84637d46032d45ad4a814597100000e7800059aa84ae891795ffff930505112d46268597300000e780c024054508c0233444012338240104ecb1a803c5150003c6050083c6250083c535002205518dc206e205d58db3e4a500b9c09104638424052d45ad4a814597100000e78040532a8aae891795ffff9305450b2d46528597300000e780001f2320040004e423382401233c4401233034032334540331a0114a631d4901154508c0e2704274a2740279e269426aa26a216182802d45ad4a814597100000e780a04daa84ae891795ffff9305a5052d46268597300000e780601923200400a9b71061833805011c65210605483e8763ee17019307f7ff10e11ce5637d1801833686ff0c622106e3f3d5fe333517011345150082800545854597100000e780601e0000411106e410610e069796ffff938646cf369610620286907588711c6e9795ffff9385b50a3d4635a8907588711c6e9795ffff9385e5082d462da021052ae01795ffff9307e5041795ffff130765053d463da0907588711c6e9795ffff9385c5012146a2604101828721052ae01795ffff9307e5fd1795ffff130705fe1d468a862e85be8597100000e780000ca2604101828082808365050005466345b60099c9054609a809466389c5000d466394c500210521a0610511a041050c6591c5086117d3ffff670023da8280397106fc22f83287ae862a8402f002ec02e802e4130500022af405659b0815822c108d472800894201460148730000006309550285456308b502914515e522751306000289456361a602130514002c001306000297300000e78080022300040009a8854511a081450ce408e805452300a400e270427421618280397106fc22f83287ae862a8402f002ec02e802e4130500022af405659b0815822c109547280089420146014873000000630b55028545630cb502914515e922751306000289456365a602130524002c001306000297300000e780e0fa01458545a300b40009a80145a300040029a081450ce408e805452300a400e270427421618280130101ba233c1144233881442334914423302145233c3143233841432334514323306143233c7141b289ae8b2a8408081306004093040040814597300000e78080e72338914005659b08c58293050141080889440146de864e8781470148730000006301950885456300b508914535ed03390141130500406372250b8545054b4a8597100000e780a0222a8aae8a0c081306004097300000e780c0ee930209c013050a402338514085659b88c58293050141130600408944de864e87814701487300000063019508630e6507114b25ed03350141094b63e8a2062330440123345401b1a8854511a081450ce408e8233004008330814503340145833481440339014483398143033a0143833a8142033b0142833b81411301014682804a85814597100000e780c018aa84ae890c084a8697300000e78000e504e0233434012338240145bf014b2334640108e823300400e3810afa528597d0ffffe78060b451bf9308d0057d558145014681460147814701487300000001a0086101a0411106e497d0ffffe78080a600008280797106f42e8813564500130f7002130710279796ffff938e66dd6363e608130f700213076102174600008338464439661b03068f05669b03b6479302c0f937e6f5051b0ef60faa86333515032d813b066502b307d600139607034992330676029355160141821376e67fbb855502be95769683471600c615c19103460600a30ff7fef69583c7150083c50500711f230fc7fea300f7002300b7007117e365defa130630066370a60493150503c99105661b06b647b385c502c5811306c0f93b86c502329546154191791f7695034615000345050093061100fa96a380c6002380a6002e85a945637cb5009305ffff130611002e961b0505032300a60005a006059305efff7695034615000345050093061100ae96a380c6002380a60093061100ae96130770020d8f1795ffff930525084285014697000000e780e000a27045618280597186f4a2f0a6eccae8cee4d2e056fc5af85ef462f066ec6ae86ee4aa8403654503ba893689328aae8b937c1500b70a110063840c00930ab00293754500ce9c89e5814b8c6085e5a1a08145630e0a005286de86038706008506132707fc134717007d16ba957df6ae9c8c6095c103bd840063ffac01218925ed83c58403054633059d41634cb60af9e1aa8c2e85c9a0807084742285a6855686de86528797000000e7806014054b0dc15a85a6700674e6644669a669066ae27a427ba27b027ce26c426da26d656182809c6c2285ca854e86a6700674e6644669a669066ae27a427ba27b027ce26c426da26d6561828780581305000383c584032ee003bc040283bd840288d8054b238c64036285ee855686de86528797000000e780e00c51f5228a33049d4105047d1451c803b60d02930500036285029665d985bf09466398c50093051500058193dc150011a0814c03bc040203bd84028458130415007d1409c803360d026285a68502966dd9054b2dbf37051100054be389a4f26285ea855686de86528797000000e780e00511fd83368d016285ca854e86829619f5b30990417d5a7d59338529016309450303360d026285a6850296050975d50da083b68d016285ca854e868296e31005ee014b23a844030265238ca402c1bd6689333b9901e1b5797106f422f026ec4ae84ee49b070600370811003a89b6842e84aa896389070114704e85b2858296aa85054591ed81cc1c6c4e85a6854a86a2700274e2644269a269456182870145a2700274e2644269a269456182805d7186e4a2e026fc4af84ef452f056ec5ae85ee483320500146933e7d2003289ae896304072a638706101c6d8146338e29018507370311009308f00d1308000f4e8601a893051600918eae962e866303640efd17adc7630fc60d8305060013f4f50fe3d105fe834516009374f40113f7f50363fa8802834526001a0793f5f503b363b7006367040383453600f614ad909a0393f5f50333e4b300458c630c64089305460055b79305260013946400598c61bf93053600b20433e4930071b7630bc6078305060063d3050493f5f50f1307000e63ede5021307000f63e9e50203471600834726001377f70393f7f70303463600f615ad9132079a075d8f1376f603598ed18d370611006386c50285c263fd2601b385d90083850500130600fc63d7c500814591e539a0e39d26ffce8599c13689ae89638b021803388500930500026372b902814e63060916ca85ce86038606008506132606fc13461600fd15b29efdf581aa13877900619b3386e940b308c90093f678008145630d3701ce87038407008507132404fc934414000506a6957df6014691ce93f788ffba9783840700850793a404fc93c41400fd162696fdf693d638009747000083b727f49744000083b224f4b714001092048504939804018508b30eb6001da013173e001a97b386c34113763e00b3f45500a181b3f55500a695b3851503c191ae9e2deaddcab6833a839305000c368e63e4b600130e000c9375ce0f139435001a94dddd81451a8745df146393c4f6ff9d8099821067c58efd8eb6959346f6ff9d82046b1982558e7d8e93c6f4ff9d829980c58e046ffd8e3696b29513c6f4ff1d829980458e7d8e13070702b295e31d87fabdb7630803029305000c63e4b3009303000c814593f633008e06106021041347f6ff1d831982598e7d8ee116b295f5f611a0814533f65500a181b3f55500b295b3851503c191ae9e63fc0e01834685030546b305d8416345d60285ce814a25a80c7508719c6dce854a86a6600664e2744279a279027ae26a426ba26b6161828709466398c600138615008581935a160019a0ae8a8145033b0502833b85020459138415007d1409c803b60b025a85a68502966dd9054a81a037051100054a638ca40283b68b015a85ce854a86829605e533095041fd597d5433058900630a350103b60b025a85a6850296050475d511a05684333a54015285a6600664e2744279a279027ae26a426ba26b61618280411106e497000000e780808f0000197186fca2f8a6f4caf0ceecd2e8d6e4dae0b2891306000232f80d46230cc10203b4090202e002e82af02ef461c003b589026307051083b409009305f5ff8e058d8113891500a10493058003330ab5026104854a17050000130b6589906001caa276027583b584ff946e829665ed08482ad803058401230ca1024c4803b509012eda033684ff0c6001ce631756019205aa95906563046601014621a08c618c61054632e02ee4033684fe833504ff01ce631756019205aa95906563046601014621a08c618c61054632e82eec0c6492052e95106508618a85029649e5c104130a8afc13048403e31b0af6b1a003ba890163080a0483b4090103b409001305faff12051181130915002104a104120a106001caa2760275833584ff946e829639e1906003b584ff8a8502960ded4104411ac104e31e0afc03b589006368a9002da0014903b589006371a90203b5090012092a99a27602758335090003368900946e829619c1054511a00145e6704674a6740679e669466aa66a066b09618280907588711c6e9785ffff9385f54f2d468287907588711c6e9785ffff9385854f39468287411106e497f0ffffe78080740000411106e497f0ffffe780a0730000757106e5014730012948bd4821a89306f6ff13d547009a92a30f56fe0507368663fcf800aa879372f50013030003e3e002ff13037005e1bf13050008198d130610086370c5021785ffff9307054e09462e85be8597000000e780e082aa60496182809305000897000000e78040560000757106e522e1a6fccaf8cef4d2f0d6ecdae8dee4e2e066fc6af86ef432892e8a014c814c81499745000003bbc5b29745000083bbc5b29745000083b4c5b200690c612ef008652aec13058a002ae01785ffff130545452ae8294d22e40da03305b6000345f5ff5915133515002300a4006265146d02758296ee8c6311051213f5f90f631b051063758901e9a8636c890d33058941b3058a014146637fc50063022c0d81463386d50003460600630da6098506e319d5fe75a013867500937686ff3386b640ad8e93b6160013371600d98ea1c20146930605ff02676297b387c5009c6313c4f7ffa58fda9733747401e18f8defb307c7009c6313c4f7ffa58fda9733747401e18f95e34106e3f9c6fc31a83387d500034707006307a7038506e319d6fe930605ffe3f9c6fa6304c5062264b386c50083c606006386a6010506e319c5fe05a0b286e296138c1600e3f026f5d29603c50600e31ba5f38149e28de28a39a04a8c8549e68dca8a63872c030345040001c96265146d11460275c265829611ed33869a41b3059a01e39a9aed0145f1bd4a8c2264f9b7014511a00545aa600a64e6744679a679067ae66a466ba66b066ce27c427da27d49618280411106e41b8605009306000802c26376d6002302b100054671a01bd6b50019ee13d665001366060c2302c10093f5f50393850508a302b1000946ada01bd6050115e613d6c5001366060e2302c10013964503699213060608a302c10093f5f503938505082303b1000d462da81396b50275921306060f2302c1001396e502699213060608a302c100139645036992130606082303c10093f5f50393850508a303b10011464c0097000000e780e0d9a26041018280397106fc907594712ae032f836f4886d906994658c612af032ec36e82ee41785ffff9305452f0a85300097000000e78080b3e27021618280086117030000670063d5411106e408611b8605009306000802c26376d6002302b100054671a01bd6b50019ee13d665001366060c2302c10093f5f50393850508a302b1000946ada01bd6050115e613d6c5001366060e2302c10013964503699213060608a302c10093f5f503938505082303b1000d462da81396b50275921306060f2302c1001396e502699213060608a302c100139645036992130606082303c10093f5f50393850508a303b10011464c0097000000e78060caa26041018280397106fc90759471986d32f836f43af0906994658c61086132ec36e82ee42ae01785ffff9305a51f0a85300097000000e780e0a3e27021618280357106ed22e926e54ae1cefcd2f8d6f42a840345050109c5833a04008544d5a0b2892e89033a840003654a03833a04009375450091e93336500163880a021785ffff9305050d35a063960a0483358a0203350a02946d9785ffff9385a50b094682961dc5814a854469a81785ffff9305850a83368a0203350a02946e05068296854441e103b689014a85d28502968da803254a038544a303910283350a0203368a022ee432e8930571022eec83250a0303068a0383360a0003378a0083370a0103388a01aaceaecc2300c10636f43af83efcc2e02800aae403b689011785ffff130545ffaae82c104a85029619e9c6652665946d9785ffff9385850109468296aa8423089400850a233054012285ea604a64aa640a69e679467aa67a0d618280397106fc22f826f44af02a841c7508719c6f3a89b684829722e8230ca10002e4a30c01002800a6854a8697000000e78060eb22658345810139c50544b9e5834591017d1513351500c264b335b0006d8d05c103c54403118901ed8c748870946d9785ffff938535f905460544829611ed8c748870946d9785ffff9385c5f1054682962a8419a03334b0002285e2704274a274027921618280411106e497f0ffffe780201600001785ffff9306a50409462e85b68517f3ffff6700634d397106fc22f826f42e848c752ae40870946d9785ffff9385a5044546829622ec2300a10202e8a30001021785ffff1306250108082c0097000000e780e0de42658345010239c50544b9e5834511027d1513351500e264b335b0006d8d05c103c54403118901ed8c748870946d9785ffff9385b5ec05460544829611ed8c748870946d9785ffff938545e5054682962a8419a03334b0002285e2704274a27421618280757106e5014730012948bd4821a89306f6ff13d547009a92a30f56fe0507368663fcf800aa879372f50013030003e3e002ff13037003e1bf13050008198d130610086370c5021785ffff930705e509462e85be8597f0ffffe780e019aa60496182809305000897000000e78040ed0000797106f422f026ec4ae84ee42a8404690865ae893309b640058d6363250308602695ce854a8697200000e780e0e0ca9404e8a2700274e2644269a269456182802285a6854a8697000000e780c0000468f9b75d7186e4a2e026fc2e966368b6042a8408659314150063639600b284a14563e39500a14493c5f4fffd9119c5106032f0054632f42af811a002f428001410268697000000e780c003a265426581cdfd55fe158505630ab50009ed97c0ffffe78060ac000008e004e4a6600664e2746161828097c0ffffe78040aa0000011106ec22e826e44ae03289aa8499cd2e84886605c18c6a91cd88624a8697c0ffffe780c0a605e180e419a023b40400854521a8630409024a85a28597c0ffffe780e0a375d1814588e423b824018ce0e2604264a264026905618280228565f5e1b703e6450308619376060189ea1376060219ea086117f3ffff6700c3ef086117f3ffff6700237b086117030000670083e3411106e422e02a8411c96347040289c9228597c0ffffe780e09e09a8054501a88545228597c0ffffe780409c19c9a285a26002644101828097c0ffffe780a09d000097c0ffffe780609c0000797106f422f026ec4ae84ee42a8904690865058d2e84636fb50283390900894533859900636cb4007d148145228697200000e780c0b8a2943385990023000500850423389900a2700274e2644269a269456182804a85a685228697000000e780e0008334090155bf5d7186e4a2e026fc2e966368b6042a8408659314150063639600b284a14563e39500a14493c5f4fffd9119c5106032f0054632f42af811a002f428001410268697000000e780c003a265426581cdfd55fe158505630ab50009ed97c0ffffe7804090000008e004e4a6600664e2746161828097c0ffffe780208e0000011106ec22e826e43284aa8499cd88660dc18c6a99cd8862228697c0ffffe780e08a19ed85458ce431a823b40400854511a88545228597c0ffffe78020887dd1814588e480e88ce0e2604264a26405618280411106e422e02a8408617d1508e005e90c70086c8c6182950870086511c5086c97c0ffffe780e084087811c5087497c0ffffe780008408647d1508e409c5a2600264410182802285a2600264410117c3ffff670003825d7186e4a2e026fc4af84ef452f056ec83ba0501368a3289aa8963e3da00d28a806108687de1286c7d5610e8637c55010870106c98651c6d4e85b2854a86d286829761a08465306463edc400b386540163ee96082c683307b600636ec7086376d70208700c6c1074147c1c6d0a85268782970345010069e9a26563e8550f286c2ce824e426866367b50eb3b6c400918c33359500558d49e5338554016363950463e7a5080c7c63eca508b3059540639745090c74a6954a85528697200000e78020a423b45901238009000868050508e8a6600664e2744279a279027ae26a616182801785ffff130505c111a81785ffff130565c029a01785ffff1305c5bff14597f0ffffe780c02f00001785ffff130595b29785ffff938685b3c1450a8689a01785ffff130585c39305f002d1bf1785ffff130595c593052003d9b7528597000000e78040a500001785ffff1305a5d69785ffff938625b89305b0021306710197f0ffffe780c04400001785ffff130545ba71b71785ffff130565bb9305e00241b7034505000e051786ffff130626df2a969786ffff938686e3369598751062146188711c6fb6858287411110650c69b29563edc50008611069fd568582637dd60028616369b502410182801785ffff1305e586a14535a01785ffff130525a99785ffff938625aae145300097f0ffffe780003c00001785ffff130535bc9305600297f0ffffe780a01f0000797106f422f0aa8502c2280050009146114497000000e78020de0345810011e942656319850203654100a2700274456182801785ffff130545c79785ffff9386c5a89305b0021306f10197f0ffffe780603500001785ffff1305f5b7b54597f0ffffe78020190000797106f422f09c6185079ce19dc7b2962ee463e6c6022a8436e83aec280097000000e78080f16265c265226608e80ce410e0a270027445618280000000001785ffff1305059f9305b00297f0ffffe780e0130000197186fca2f8a6f4caf0ceecd2e8d6e4dae05efc03bb050003370b00846594692a89130517002330ab006dcd5ae409072330eb0065cbb28a36f85af02e8597000000e78060f09385440063ef950caa892ef4081097000000e78000ef8d4563faa50c09811304f5ff63fe8a02938b1a0013952b0026956364950c2af4081097000000e78060ec2a8a63998b0233854401636c950a2ae863f649051785ffff13050594f1a015452304a900233009005a8597000000e78020c3b1a08a0a33859a002105636895082af4081097000000e780a0e7b385440163e39508aa892ee863644509338549412aec280097000000e78080df6265c26522662338a9002334b9002330c9005a8597000000e780c0bde6704674a6740679e669466aa66a066be27b09618280000000001785ffff1305258b3da81785ffff1305259fb9451da81785ffff1305c58925a01785ffff1305258939a81785ffff1305858811a81785ffff1305e58729a01785ffff130545879305b00297f0ffffe78020fc0000397106fc22f826f42a8402e408083000a146a144a28597000000e78060ba0345010105e16265631f9502a264086097000000e78080b32685e2704274a274216182801785ffff1305c5a29785ffff938645849305b0021306710297f0ffffe780e01000001785ffff13052595b94597f0ffffe780a0f40000397106fc22f826f42a84a307010008081306f10085468544a28597000000e780a0b2034501010de16265631095048304f100086097000000e780a0ab2685e2704274a274216182801785ffff1305e59a9775ffff9386657c9305b0021306710297f0ffffe780000900001785ffff1305258eb54597f0ffffe780c0ec00005d7186e4a2e026fc4af8ae842a898c69054632e002e402e889c90a8597000000e780e0910266426411a001442808a685a28697000000e78040a9034581011de5027563168504c2652266826688602338b9002334c9002330d900a6600664e27442796161170300006700c3a01785ffff1305c5909775ffff938645729305b0021306f10297f0ffffe780e0fe00001785ffff1305d584c94597f0ffffe780a0e20000011106ec22e826e49c692a84637df700b384e74063e3d400b684b306970063ede60263f7d7001545a300a400054531a8998e639dd4028c61ba953285268697100000e780204e014504e42300a400e2604264a264056182801775ffff1305e56bf14597f0ffffe780e0db00002685b68597f0ffffe780605400005d7186e4a2e026fc4af84ef452f02e8483b905012a896145a14597b0ffffe780001a59c1aa84086888e8086488e4086088e0054a52e402e802ec1314ba002800a28597f0ffffe780c07d13050006a14597b0ffffe780a01621c923304501233445012338050004ed9775ffff9385c5760cf1a2650cf5c2650cf9e2650cfd23303505233405042338050420ed23340900233839012330a900a6600664e2744279a279027a6161828097b0ffffe780201300000c6591c5086117b3ffff6700a31082805d7186e4a2e026fc4af8ae84806590612a892800a28597e0ffffe780c03c0345810019c5426529e109452300a90029a805040dc09305910080e4130610024a8597100000e780403aa6600664e2744279616182801775ffff13056572f14597f0ffffe78060c8000097e0ffffe78080570000357106ed22e926e54ae1cefcd2f8d6f4daf02e89aa8a2800d68597000000e78040f7034581008944630b951675cd0345210283451102034631028346410222054d8d4206e206558e518d83456102034651028346710203478102a205d18dc2066207d98ed58d82154d8daae40345a101834591010346b1018346c10122054d8d4206e206558e518d8345e1010346d1018346f10103470102a205d18dc2066207d98ed58d82154d8daae00345210183451101034631018346410122054d8d4206e206558e518d83456101034651018346710103478101a205d18dc2066207d98ed58d82154d8d2afc0345a100834591000346b1008346c10022054d8d4206e206558e518d8345e1000346d1008346f10003470101a205d18dc2066207d98ed58d82154d8d2af829a082e482e002fc02f803b58a010c6903b40a0113060002639bc5040c6108181306000297100000e78000650125854421e103b50a0210610818a28597e0ffffe7800029c279638f09120665627bc145637fb50263070b004e8597b0ffffe780e0f08144130550032300a90011a08544050475c823b88a002685ea604a64aa640a69e679467aa67a067b0d6182804145814597f0ffffe780604e2a892e8a4146ce8597100000e780a01a0345190083450900034629008346390022054d8d4206e206558e518d83455900034649008346690003477900a205d18dc2066207d98ed58d8215c98d03459900034689008346a9000347b9002205518dc2066207d98e0346d90033e7a6000345c9008346e90022068347f900498ec20603b58a02e207dd8e558e14651c610216598e3696be9533b7f5003a966304d6003337d60015ef0ce110e563070a004a8597b0ffffe780e0e163070b004e8597b0ffffe78000e103b40a0131b71775ffff1305c547f14597f0ffffe780c09d00001775ffff13058546f5b71775ffff1305e5479775ffff9386654a9305b002900897f0ffffe78020b600000e059775ffff938545c82e950c6105458285094582800d4582801145828097e0ffffe78060280000357106ed22e926e54ae1cefcd2f8d6f4daf02e8a2a8908100546814597e0ffffe7802006034501020dc12275c27597000000e780a0faea604a64aa640a69e679467aa67a067b0d61828003156102831541020356210283461102231ea104c205d18da274627503560104c27aaeccaae42318c104f5c603150105a6652314a1002ee013050002130b0002814597f0ffffe78000322a84ae89ac08194697100000e780204313d58403a306a40013d504032306a40013d58402a305a40013d504022305a40013d58401a304a40013d504012304a40013d58400a303a4002303940013d58a03a30aa40013d50a03230aa40013d58a02a309a40013d50a022309a40013d58a01a308a40013d50a012308a40013d58a00a307a40023075401130564018a85294697100000e780c0f58144631c6a01130600022285ca8597100000e780e0369334150063870900228597b0ffffe78000c513057004e38f04ec0145e1bd3945d1bd130101c0233c113e2338813e2334913e2330213f233c313d2338413d2334513d2330613d233c713b930700026312f6523a8ab6892a8903c5950103c6850183c6a50103c7b5012205518dc2066207d98e558d03c6d50183c6c50103c7e50183c7f5012206558e4207e2075d8f598e0216518d2af003c5150103c6050183c6250103c735012205518dc2066207d98e558d03c6550183c6450103c7650183c775012206558e4207e2075d8f598e0216518d2aec03c5950003c6850083c6a50003c7b5002205518dc2066207d98e558d03c6d50083c6c50003c7e50083c7f5002206558e4207e2075d8f598e0216518d2ae803c5150003c6050083c6250003c735002205518dc2066207d98e558d03c6550083c6450003c7650083c575002206558e4207e205d98dd18d82154d8d2ae413050002854597b0ffffe780c0af630505402a8413060002814597100000e78060d01145854597b0ffffe780c0ad6305053eaa84a301050023010500a30005002300050013050002930b0002814597f0ffffe780c00c2a8bae8a2c001306000297100000e780e0d8228597b0ffffe78000aa13054a0063634537814597f0ffffe780e009aae2aee682ea2320412dd00588028c0597f0ffffe78060f2338649018802ce8597f0ffffe78060f1166ab6695664268597b0ffffe78060a5dae2d6e6deead2eecef2a2f68945130514032308b116636a8530814597f0ffffe7802004aae4aee882ec0d4597e0ffffe780a0832330a12c2334b12c2338012c99c1814511a8880597e0ffffe78080908335012d0335012c8e052e95c1450ce18335012dd6698505138409012338b12c6362342d0335812c6399a500880597e0ffffe780208d8335012d033a012c13953500529500e19384150005042338912c630f04280335812c639ca4008805a68597e0ffffe780008a8334012d033a012c939a340033055a0100e136752295636d85262ad47010a8002c1097f0ffffe78040e2033b812c7d556384a4026410a10a52850c61130485002ed4a8002c10268697f0ffffe780e0dfe11a2285e3930afe63070b00528597b0ffffe78080939665801a33863501a80097f0ffffe78060dd13061117a800a28597f0ffffe78060dcf66536762e96a80097f0ffffe78060dba669c66a3665666a11c5166597b0ffffe780208f167511c5766597b0ffffe780408e82e002fc02f802f40403c802801a1306c002814597100000e780e0ad130680132685814597100000e780e0ac1775ffff9305b5cb4146228597100000e78080b8370501011b0505022320a114233c012a88051306800f814597100000e780a0a988058c0297b0ffffe780a0baa8008c051306800f97100000e780c0b4a800ce85528697b0ffffe78060c28802ac001306800f97100000e780e0b2880513060004814597100000e78000a5033581229305000263eaa50a5a655de5033501229a653386a50032e3ba66b335b600b6952ee78345012399c1fd552eeffd55130610082eeb6379c5121306000800136309c500098e2295814597100000e780c09f88028402a28597b0ffffe78000c821459305312c9060a38ec5fe93568600238fd5fe93560601a38fd5fe935686012380d50093560602a380d500935686022381d50093560603a381d50061922382c5007d15a104a1055dfd0336812228108c0597100000e78020a62c10130600024a8597100000e78020a563870a004e8597a0ffffe78000768330813f0334013f8334813e0339013e8339813d033a013d833a813c033b013c833b813b1301014082801775ffff1305858925a01775ffff1305e58839a81775ffff1305458811a81775ffff1305a58729a01775ffff13050587f14597e0ffffe780002e000097a0ffffe780a07000001775ffff130525d89775ffff9386a5dc9305b002900297e0ffffe780604600009305000897f0ffffe780e0a30000697106f622f226ee4aea4ee652e2d6fddaf9def5e2f1e6ed2e8a2a89014481490d45aae082e49304110501163335c00093b51500b36ab500130b1108894b7d5c88088c0097f0ffffe7806057034501056309751f6301051003c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8d2ae903c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8d2ae503c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8d2ae103c5140083c5040003c6240083c6340022054d8d4206e206558e518d83c5540003c6440083c6640003c77400a205d18dc2066207d98ed58d82154d8daafc63890a00dda002e902e502e182fc639e0a0ca81813060002d28597100000e780c0c5012579e1639a091628110d46a28597e0ffffe780e0892a7559c96a75ca752a76aae9aee5b2e1a8188c0197f0ffffe780c0350305eb008305db000346cb00e6792303a10aa205d18d2312b10a03459b0083458b000346ab008306bb0022054d8d4206e206558e518d2ad103451b0083450b0003462b0083463b0022054d8d4206e20683455b00558e518d03464b00a20583466b0003477b00d18d834c0108c2066207d98ed58d82154d8d2aed11a081496a658a550316410a8306610a2af82edc231ec102230fd102630e8409050401b5638609060305e1038315c1036256c2762307a1022316b10232d436f0130511010c103d4697000000e78080734ee423089101a8182c00054697f0ffffe78000ef667535c92a658a656676aaf0aeecb2e8880897f0ffffe78020052334a9004e8597f0ffffe780a0ba014531a01305a005a300a90005452300a900b2701274f2645269b269126aee7a4e7bae7b0e7cee6c556182801775ffff1305e5a5f14597e0ffffe780e0fb00001775ffff1305a5ad9305b002edb71775ffff1305c5a59765ffff9386c5309305b002900897e0ffffe78000140000717106f522f126ed2a8432e402ec02e802fc02f8a303010232f4aee02800aae40808aae813057102aaec28109305710297f0ffffe780402e058901e9034571020dc9a300a40005450da888102c101306800397000000e7804063f954ca65881097f0ffffe780402b058969d991ccfd14f5b7c26562660ce810ec2300a400aa700a74ea644d61828097a0ffffe780c03300004d7186e6a2e226fe4afa4ef652f256ee5aea5ee662e2e6fdeaf9eef5b2842e8a2ae0014c814d8149814b1304110cfd5a3d4d32e82ee48801e285268697d0ffffe780c0530345010c631e052863045c3103459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8d2ae90345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8d2ae503459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8d2ae10345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8daafca81813060002d28597100000e780c08c0125631305188801e285268697d0ffffe78000510e6b630d0b1ece6c2e65637f9d15aaeceef04145814597e0ffffe780e079aa84ae8b4146da8597000000e780204683c5840083c9940003caa40083cdb40003c6c40003cdd40083c7e40083caf40003c3040003c7140003ce240083c6340003c8440083c3540083c8640083c2740063870b04268542f4c68496e01a896af01e8d52ec728a6ef8b68dcee4ba89b2e856fcbe8aae8b97a0ffffe7800011de85d687e27a46664e87a669ee86c27d528e626aea83027d4a838662a68822780675631f0514a20933e5b900420ae20db3e54d014d8d220db365cd0013960701e20a33e6ca00d18d821533e9a500131587003365650093150e0113968601d18d4d8d93958300b3e505011396080193968201558ed18d82154d8daaf093840cff130a0b012685814597e0ffffe7800069aa8cae8bd285268697000000e7804035e6e1dee5a6e928118c0197f0ffffe780c0e90c1988618c65814baa7daaf4aef88549c264226afd5a3d4d666511c55a8597a0ffffe7808003050c91bb2e6586765de533e5790111cd638c0d024675a675026608f20cee14e2233426012338b6013da01305500382652380a50023b80500638f0d006e8597e0ffffe780407801a81305200382652380a50023b80500b6601664f2745279b279127af26a526bb26b126cee7c4e7dae7d716182801765ffff13056563f14597e0ffffe78060b900001765ffff130525649765ffff9386a5669305b002301197e0ffffe78060d200001765ffff1305d56b93059002e9b797d0ffffe780a0450000757106e522e1a6fccaf8cef4d2f02a89814432e402e81304910181153335b00093351900b369b500094a28082c0097f0ffffe78020e40345810165d9630c451303459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8daaec0345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8daae803459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8daae40345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8daae0e39909ee880013060002ca8597000000e78080530125e31e05ec93f4f40f850413f5f40fe30795ec1765ffff1305a548f14597e0ffffe780a09e00002685aa600a64e6744679a679067a4961828071c693f7f50f2300f5003307c500a30ff7fe894663fcc60aa300f5002301f500230ff7fea30ef7fe994663f1c60aa301f500230ef7fea14663fac60893f5f50f9b9785003307a0400d8bad9f198e9b950701ad9f2a97719a1cc3b305c70023aef5fe63f5c6065cc31cc723aaf5fe23acf5fee14663fcc604137847005cc71ccb5ccb1ccf6108939807029396070293d8080223a2f5fe23a4f5fe23a6f5fe23a8f5fe33060641fd474297c69663f0c7020116937706fe93870702ba9714e314e714eb14ef13070702e31af7fe8280397122fc26f84af44ef052ec56e85ae45ee093f735006387074069c2aa8719a06303062a83c60500850513f735002380d7007d1685076df793f637003e87cdea3d48637dc804930806ff6378180133e8b700137878006304083093d84800138f1800120f2e9f2e87be86832e0700032e4700032387000328c70023a0d60123a2c60123a4660023a606014107c106e31eeffc85089208c695c6973d8a137886001377460093762600058a630c080083a8050003a84500a107a10523ac17ff23ae07ff11c798419107910523aee7fe6391061e09c603c705002380e7006274c27422798279626ac26a226b826b216182807d476379c70a094883c805009841638806290d486386061d9306c6fe03c3150003c8250093f306ff13843700938435009382330123801701a38067002381070113d94600ae92a687a28803a8170083a5570083a697001b53870103a7d7009b1f88001b9f85009b9e86001b5888019bd585019bd686011b1e87003363f3013368e801b3e5d501b3e6c60123a0680023a2080123a4b80023a6d800c107c108e39657fa9307190092073516b385f40033067640a29793780601137886009376460013772600058a6384080883cb050003cb150083ca250003ca350083c9450003c9550083c4650003c4750083c3850083c2950083cfa50003cfb50083cec50003ced50003c3e50083c8f50023807701a380670123815701a381470123823701a382270123839700a383870023847700a38457002385f701a385e7012386d701a386c70123876700a3871701c105c1076304080483c2050083cf150003cf250083ce350003ce450003c3550083c8650003c8750023805700a380f7012381e701a381d7012382c701a382670023831701a3830701a105a1079dc203c3050083c8150003c8250083c6350023806700a380170123810701a381d70091059107e30307e283c6050003c715008907238fd7fea38fe7fe890539b513f73700e31d07ec39b59306c6fe93f306ff1384170093841500938213012380170113d94600ae92a687a28803a8370083a5770083a6b7001b53870003a7f7009b1f88011b9f85019b9e86011b5888009bd585009bd686001b1e87013363f3013368e801b3e5d501b3e6c60123a0680023a2080123a4b80023a6d800c107c108e39657fa9307190092073d16b385f40033067640a297a1b593d84800938e18002e88033e88000333080085062334c7012330670041084107e3e5d6ff85089208c695c6973d8a01bb9306c6fe03c8150093f306ff13842700938425009382230123801701a380070113d94600ae92a687a28803a8270083a5670083a6a7001b53070103a7e7009b1f08011b9f05019b9e06011b5808019bd505019bd606011b1e07013363f3013368e801b3e5d501b3e6c60123a0680023a2080123a4b80023a6d800c107c108e39657fa9307190092073916b385f40033067640a29749b3aa8709b919ca0347050083c705007d166317f700050585057df6014582800345050083c705001d9d8280aa862e87b287630db50cb388c5403308c040b388a84006082e832a8e6372181b3346b5001d8a637fb50a63010612cdcb1386f7ff9d4563f8c51813061700b305c54093b5750093c5150093f5f50f638a0516b365e5009d896395051693f587ffba95033603002103210e233ccefee39a65fe13f687ff13f57700aa87b385c600329739cd0345070005462380a5006389c704034517000946a380a5006382c704034527000d462381a500638bc702034537001146a381a5006384c7020345470015462382a500638dc700034557001946a382a5006386c700834767002383f5003685828029ea3306f5001d8a65ca1386f7fffdd7b307c5007d5821a07d16e30106ffb305c70003c5050093f57700fd17a380a700e5f59d4763fac70ab2871d48e117b305f7008861b385f60088e1e369f8fe93777600cdd7fd173306f700834506003386f6002300b600f5b71376750041ca9385f7ffc9d72a867d5821a0fd15e38005f903450700050693777600a30fa6fe0507edf79d4763fcb704938885ff93f888ffa10833051601ba8703b807002106a107233c06ffe31aa6fe469793f77500130617008ddfba9711a005060347f6ff0505a30fe5fee31af6fe36858280cdba3685d5b713061700f9bfb287a5b73285ae8713061700e1f919b73e8625bf2a86be8549bf0000d182e6ad7f520e5108c9bcf367e6096a1f6c3e2b8c68059b3ba7ca8485ae67bb6bbd41fbabd9831f2bf894fe72f36e3c79217e1319cde05bf1361d5f3af54fa54b598638d6c56d340101010101010101ff00ff00ff00ff00fffefefefefefefe80808080808080800a0a0a0a0a0a0a0a0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008cd0900000000000010000000000000040000000000000008bd01000000000000100800000000004000000000000000010000000000000060090100000000000000000000000000011101250e1305030e10171b0eb44219110112060000023901030e0000032e001101120640186e0e030e3a0b3b053f198701190000041101250e1305030e10171b0eb44219110155170000052e006e0e030e3a0b3b05200b0000062e001101120640186e0e030e3a0b3b050000072e006e0e030e3a0b3b0b200b0000082e011101120640186e0e030e3a0b3b0b360b0000091d00311311011206580b590b570b00000a1d0031135517580b590b570b00000b1d00311311011206580b5905570b00000c1d0031135517580b5905570b00000d2e006e0e030e3a0b3b0b3f19200b00000e2e011101120640186e0e030e3a0b3b0b3f1900000f1d0131135517580b590b570b0000101d01311311011206580b590b570b0000111d01311311011206580b5905570b0000121d0131135517580b5905570b0000132e006e0e030e3a0b3b053f19200b0000142e011101120640186e0e030e3a0b3b05360b3f190000152e011101120640186e0e030e3a0b3b053f190000162e0111011206401831130000172e0011011206401831130000182e001101120640186e0e030e3a0b3b0b0000192e011101120640186e0e030e3a0b3b0b00001a2e011101120640186e0e030e3a0b3b0500001b2e001101120640186e0e030e3a0b3b0b3f1987011900001c2e006e0e030e3a0b3b0b870119200b00001d2e011101120640186e0e030e3a0b3b05360b3f198701190000004d0000000400000000000801962900001c00d4420000000000002c120000e8420100000000000e00000002452d0000020000000003e8420100000000000e0000000152914b000064350000010b02000000c62200000400000000000804962900001c00201600005c0000002c1200000000000000000000700e00000201190000021f050000057d0c00005616000002f9050106b477010000000000020000000152dc3200002b0c000002eb0102323c0000029730000005e6350000982300000693030105e6350000982300000693030105e6350000982300000693030105e6350000982300000693030105e6350000982300000693030105c5280000ec21000006930301050c2b0000dc4500000693030105573800006f3700000693030105c50b0000f90300000636050105e63500009823000006930301000002ad0c0000029730000005353f0000982300000801040105353f0000982300000801040105353f0000982300000801040105353f0000982300000801040105353f0000982300000801040105b03000005317000008010401054d0b0000d534000008010401000005a6000000844600000273040105fe120000de40000002730401052f4500002b050000024905010506080000cc000000024905010536280000f903000002610601000293300000025c120000029031000007124800007527000003d0010002023e00000737130000d3450000038e01072c3b000093300000038901072c3b00009330000003890100000269480000028a2e000008b677010000000000420100000152c21500007635000005d303096500000026780100000000000200000005f1360a2c1900000000000005f115097200000038780100000000000200000005f2360a391900004000000005f215097f00000080780100000000000200000005fd360a461900007000000005fd1509f30000008e780100000000000200000005fd470b00010000a878010000000000020000000503011e0b8c000000ba7801000000000002000000050701360c53190000a0000000050701150b0d010000c87801000000000002000000050701470b1a010000d67801000000000006000000050f0133000002a30b000007682b00005d3b000005430107e52d00006f29000005430100024b2900000d02140000d81b00000587010002ff4300000dd0460000ba380000052a010002771400000e76800100000000007000000001522a2e000093300000059a0fd902000020090000059b1110a21a00007c8001000000000008000000054e1d110d1a00007c80010000000000080000001af8020909410100007c80010000000000080000001cef5000000af70200005009000005511c09201f00008e800100000000000400000005511609090300009c80010000000000080000000551280f942100008009000005651412571b0000b0090000225901090a441b0000e0090000181209000000000002650700000d73320000d81b000005870100026f0700000e06870100000000007000000001521f03000093300000059a0fe5020000800d0000059b1110f61a00000c8701000000000008000000054e1d110d1a00000c87010000000000080000001af8020909410100000c87010000000000080000001cef5000000ae2030000b00d000005511c092d1f00001e870100000000000400000005511609090300002c87010000000000080000000551280fa1210000e00d000005651412631b0000100e0000225901090a441b0000400e000018120900000000000002ec49000013370a00006c0a000009bd0601137f0300008e2e000009f6060113de480000ca4000000910070105b90c000023050000096e050114f878010000000000e4010000015289020000cc31000009de04030bbc04000016790100000000000c00000009e504130bc904000032790100000000000400000009ea04190bd60400006e7901000000000002000000090a051a12e3040000d00000000917052411131d0000567a010000000000040000000980051211001d0000567a010000000000040000000fc702090b4c1f0000567a010000000000020000000f6d020c000000127511000010010000091a051112201d0000400100000994041212001d0000700100000fc702090c4c1f0000a00100000f6d020c00000012fc1e0000d0010000090b05200b50010000e87901000000000006000000149403160b6a010000fc7901000000000004000000149503090012091f000000020000090c05210b5d010000ee7901000000000004000000149403160b77010000007a01000000000004000000149503090011e30400001a7a0100000000001a000000090e052411131d0000207a010000000000040000000980051211001d0000207a010000000000040000000fc702090b4c1f0000207a010000000000040000000f6d020c00000011b81d000044790100000000001c00000009eb041610531d000044790100000000001c00000013310910471d000044790100000000001c00000012200910ab1c000044790100000000001c00000012874c101e1c000044790100000000001c00000011533111511c000044790100000000001c0000000b940d0910811c000044790100000000001c0000000d321110111c000044790100000000001c000000107c091270190000300200000bb0091d10b21900005079010000000000020000000a2b3509270100005079010000000000020000000a5352000012931c0000800200000bb1091510c11c000052790100000000000800000010541c10641d0000527901000000000008000000115016090f1e000052790100000000000800000012871f000009621c00005c79010000000000020000001054150000000000000000000015327b0100000000007803000001528d470000202e0000093c0512c01f0000b0020000093e05170cb31f0000e00200001583020f00116a1e0000607b0100000000000400000009470525115d1e0000607b010000000000040000001741033311201a0000607b010000000000040000001708032711be190000607b010000000000040000001ae502090999000000607b010000000000040000001c62500000000011381c0000647b010000000000da00000009470523112b1c0000647b0100000000006e0000000b8b010912d61d0000100300000b5801100fc41d000040030000138c190f1b1e000070030000132c120970190000887b010000000000040000000c260e09331e0000a07b010000000000040000000c3212093f1e0000ac7b0100000000000a0000000c3913094b1e0000c27b0100000000000a0000000c412509271e00009c7b010000000000040000000c2e10000000112d1d0000847b010000000000040000000b57011211001d0000847b010000000000040000000fc702090b4c1f0000847b010000000000020000000f6d020c00000011d61d0000f07b0100000000004e0000000b8c010910c41d0000f07b0100000000004a000000138c19101b1e0000f07b0100000000004a000000132c120970190000f07b010000000000040000000c260e094b1e0000287c0100000000000c0000000c4125093f1e00001c7c010000000000040000000c391309331e0000187c010000000000040000000c32120000000012831e0000a0030000094c051312a81e0000d003000017b9010911771e00003e7c010000000000120000001914010c102d1a0000447c0100000000000400000017dc1f0b0e1b0000447c010000000000040000001a5a010f000000000ccd1f000000040000094c051c11b81d0000727c010000000000720100000959052310531d0000727c0100000000007201000013310910471d0000787c0100000000001e00000012200910ab1c0000787c0100000000001e00000012874c101e1c0000787c0100000000001e00000011533111511c0000787c0100000000001e0000000b940d0910811c0000787c0100000000001e0000000d321110111c0000787c0100000000001e000000107c091270190000300400000bb0091d10b2190000847c010000000000020000000a2b350927010000847c010000000000020000000a5352000012931c0000800400000bb1091510c11c0000867c0100000000000800000010541c10641d0000867c01000000000008000000115016090f1e0000867c0100000000000800000012871f000009621c0000907c010000000000020000001054150000000000000010711d0000967c0100000000004e010000122209103a1a0000967c01000000000014000000123a270b84010000967c010000000000060000001ad60d1f11541a00009c7c010000000000080000001ada0d200b471a00009c7c010000000000080000001a460617000b611a0000a47c010000000000060000001adb0d240010471d0000aa7c0100000000001a00000012471510ab1c0000aa7c0100000000001a00000012874c101e1c0000aa7c0100000000001a00000011533111511c0000aa7c0100000000001a0000000b940d0910811c0000aa7c0100000000001a0000000d321110111c0000aa7c0100000000001a000000107c091270190000b00400000bb0091d10b2190000b47c010000000000020000000a2b350927010000b47c010000000000020000000a5352000012931c0000000500000bb1091510c11c0000b67c0100000000000800000010541c10641d0000b67c01000000000008000000115016090f1e0000b67c0100000000000800000012871f000009621c0000c07c010000000000020000001054150000000000000010471d0000c67c0100000000001c00000012473510ab1c0000c67c0100000000001c00000012874c101e1c0000c67c0100000000001c00000011533111511c0000c67c0100000000001c0000000b940d0910811c0000c67c0100000000001c0000000d321110111c0000c67c0100000000001c000000107c091270190000300500000bb0091d10b2190000d27c010000000000020000000a2b350927010000d27c010000000000020000000a5352000012931c0000800500000bb1091510c11c0000d47c0100000000000800000010541c10641d0000d47c01000000000008000000115016090f1e0000d47c0100000000000800000012871f000009621c0000de7c0100000000000200000010541500000000000000107d1d0000187d01000000000012000000125a120939200000247d01000000000004000000127f0e0010fb190000467d01000000000006000000125019107b1a0000467d010000000000060000001c1a0e11ca190000467d010000000000060000001ae5020909a6000000467d010000000000060000001c62500000000a7c190000b00500001250190a891d0000f005000012541b0f881900006006000012631a10d6190000b87d010000000000020000000a2b350934010000b87d010000000000020000000a5352000009951d0000ba7d0100000000000c00000012641b10a11d0000d07d010000000000120000001266160946200000dc7d01000000000004000000127f0e00096e1a0000427d01000000000004000000124f2c10e81900002e7d01000000000010000000124a12119b1f00003a7d010000000000040000001ccb051b118d1f00003a7d010000000000040000000e7e04080b7b1f00003a7d010000000000040000000e2e030900000000000012e3040000b00600000963052811131d0000407e010000000000040000000980051211001d0000407e010000000000040000000fc702090b4c1f0000407e010000000000020000000f6d020c00000011751100006c7e010000000000260000000965051512201d0000f00600000994041212001d0000200700000fc702090c4c1f0000500700000f6d020c000000000d28380000d52d000009f201135e1700005e2b000009f4050113123100003e2900000943070105412700006a1c0000099c040116a8850100000000009800000001526211000011f9160000b4850100000000001800000009e6071b0b65100000b4850100000000000c0000001f1701120011c1160000da850100000000005800000009e807091168210000e4850100000000004a0000001f65012711b5150000e685010000000000480000002027051611c9150000fa85010000000000060000001f66013c0bc9040000fa85010000000000060000001f700109000b651000000286010000000000140000001f6701150b651000001886010000000000160000001f69011100000000131f0700007e23000009e507010002451a0000051f170000222f0000099304010002282f000002cc31000006dc7a0100000000005600000001529c490000ff19000009f304000005fa080000584900000964040105420f00001f0900000979040115b87e0100000000007e010000015231390000222f00000938040c59100000800700000939041912db1c0000b0070000094d041d0a94190000e00700001d2f110012a9110000100800000956041a11b6110000407f01000000000018000000096b04150bb3010000467f010000000000120000000981042c0011b6110000667f01000000000018000000096c04190bb30100006c7f010000000000120000000981042c0011881a0000867f010000000000040000000973041f111a1b0000867f010000000000040000001a96011a09b3000000867f0100000000000400000018ee1c00000bbf0100008a7f010000000000080000000976040b0012e71c000040080000093f041d0aa0190000700800001d2f11000bcb010000d87f0100000000000a0000000946041512951a0000a0080000095d042612261b0000e00800001a5a010f10321b000006800100000000000400000018d93609c000000006800100000000000400000018ee1c0000000002f101000007ab3c0000a93800001f550102d83700000ee680010000000000bc01000001527e3500005e2b00001f1f0ffb1d0000100a00001f201212e81d0000400a0000133f050911e71e00006c81010000000000d40000001372020f11bc1a0000768101000000000008000000249e01320b751b00007681010000000000080000001a5a01090011bf1b00007e81010000000000ac00000024a2012209cb1b000084810100000000001a000000252c1010d71b00009e810100000000008c000000252f0510cd0000009e810100000000000c0000002552160b840100009e810100000000000c000000064005160010ef1b0000e4810100000000000a000000256a160960200000e481010000000000020000002514070010e31b0000ce810100000000000a0000002569160953200000ce81010000000000020000002514070009da000000c2810100000000000400000025651b09cb1b000016820100000000001400000025771609cb1b0000f68101000000000012000000255a1e000011c91a000036820100000000000200000024b701430b751b00003682010000000000020000001a5a010900116c1f000038820100000000000400000024b8011c11ac1b00003882010000000000040000000ea9050d098e1b0000388201000000000004000000231a0900000000000f901e0000700a00001f252712d41e0000a00a0000175f040d12c11e0000d00a00002445022912af1a0000000b000024de0309115f1f000048810100000000000a0000001a09091311a01b000048810100000000000a0000000ea9050d098e1b000048810100000000000a000000231a09000000000000000002383d000002b94400000592040000752700001f3501010002f81900000523230000752700001f65010100000264290000055c490000714600001f6f0101158884010000000000200100000152bd090000b94400001f3401125b210000b00b00001f35012311a2150000ac84010000000000de0000002027051612c9150000e00b00001f3601100cc9040000100c00001f700109000b65100000d484010000000000160000001f3801150c65100000400c00001f4101110b7b2100000a85010000000000020000001f41011112d4160000700c00001f3c01220f7f100000b00c00001f1a0911eb1600002a850100000000000a00000009a3041209da1f00002a850100000000000a0000001f1a260000000b651000007685010000000000120000001f3e011100000013e41c0000f81900001f63010100027847000007a91c0000e02d00001f15010002f108000002e02d0000070b350000752700001f1a0100000555310000132300001f13010100020f30000016a282010000000000b400000001526b17000010b8220000b0820100000000009600000009a41a11a6220000b082010000000000960000002679022a0c99220000300b000026b6060f0000001756830100000000003800000001527717000007741800001530000009a3010788440000664b000009bf01000297300000188e830100000000000a0000000152bc470000eb41000009c6199883010000000000b60000000152164200001530000009ca106b170000a683010000000000a200000009cb0910b8220000a8830100000000009600000009a41a11a6220000a883010000000000960000002679022a0c99220000700b000026b6060f00000000194e840100000000003a000000015282370000664b000009ce09771700006e840100000000001400000009cf090000027809000005db0f00009330000009bb09010002210c00001a4e860100000000001600000001524b3000002610000009d0080b3d1800004e860100000000001600000009d0083e000000027839000002e3490000026248000019a27701000000000004000000015282090000ca4b000001fa10a1010000a2770100000000000400000001fa050934000000a2770100000000000200000003d21e000000000002812700001ba6770100000000000e00000001521d0e00008347000004341baa7e0100000000000e0000000152f3150000242e0000046e1ce73c00000a1200000495011c6c0f00004b31000004850100027c39000005f90900008f100000075f0a0105f90900008f100000075f0a0105f90900008f100000075f0a0105f90900008f100000075f0a0100029d31000002211d000002a02300000766330000194500000a7c0107b23a0000c10100000a7c0107922a0000fd4000000a7c0107804a0000e13d00000a7c0107201b00008d3c00000a7c010002383600000712000000241a00000a4b0107522d00001e4900001c5b0107e1310000fc2100001c5b01070c2200004b3400000a4b010002764a000005ef360000fd4000001cc7050100029730000007c20a00009c3a00001c190100029b0b0000079a1b0000b34100001cd90100000297300000058b110000511a00001ae4020105d01a0000272800001a56010105b4430000a54600001acb0d0105ac250000823d00001a98060105b3050000993d00001a4206010519410000b00800001a860d010565280000b12800001a16040105e13700008b3a00001ae40201057a190000d21100001a8f0101056d4100006a2f00001a5601010546260000280900001af7020105a90d0000f11700001a040901054c040000d01900001a560101054c040000d01900001a560101020f0700000340860100000000000e00000001526e420000663900001a0b0d000546260000280900001af702010002b403000002d8370000074a050000d931000018d70107613400001729000018e30107400d00000012000018d701070b3e0000fe30000018e30100027937000005fa010000f945000018ec0101000297300000077b2f000093170000181101077b2f0000931700001811010002383d000005ea140000d9310000185f0101000002ec0c000002264900000781140000843b000023520100029730000007de1b00002d3d000023190107de1b00002d3d0000231901000002d92d000007ff170000d92d000025290107923b0000ca3b00002534010d374700005b1c0000254701079d0f00007f3e0000251301079d0f00007f3e0000251301000002211d0000024b2d000002d7290000020c430000055f120000ab2300000baa0901053c3c0000833f00000b8f0d01057b360000f60000000b560101053a080000e10e00000b8a0101000002a710000002ad100000078b270000873900000d310102b50c00000756400000b71000000d350100000000027b46000002982e000002d8370000079c2e0000261d00001078010002fd4900000721430000431f0000105401000002f649000002d837000007790700009f120000114d01020c0000000222450000076b160000590000001150010000000002161b000002f108000007fe050000022600001d2e01076d130000532200001d2e01000000022d08000002d83700000556450000f12000000f6c020100028f4600000502210000fd4000000fc602010502210000fd4000000fc602010502210000fd4000000fc602010000000208000000020c0000000d760a00000c1a0000128601074e0e000015430000121a01020c1a000007e51e000075270000128701000d790800006b19000012260107a63d000024130000127a01074b2a0000d2010000127201074b2a0000d201000012720107a63d000024130000127a010002211d00000297300000076d4800000c00000013300107064a00001f010000132901000226490000075a1a00001f010000138a010002f62f00000597260000b00b0000136c02010002e141000005092c000004300000133e0501000002b60a000007413d00007b3c00000c180107e0290000c23600000c240107030f00001f2a00000c0b010797210000d92100000c11010797210000d92100000c11010797210000d92100000c1101000297300000053d360000e33300001707030105e1270000984600001740030107f60c00002f2a000017d30105e93300002534000017b80101050a0400001d3d0000175b040100024b2d000002a73000000524010000460500001913010100000222470000024b29000005fa4a00002a47000024dd030100028f46000005e52600002a47000024410201000297300000058b2c000026320000249b0101000000022b45000005533a0000371a0000148f030105a3310000820e0000148f030102a32b0000026b1400000531440000c646000021e801010531440000c646000021e8010100000002ec0c000002f00c000002ec0000000506190000e03300000e53050100020a23000005c0380000552900000ea8050105c0380000552900000ea8050100000509440000312f00000e930401026b370000052f490000402a00000e2a03010005cc080000402a00000e7d040100023308000002a030000005a40e0000370500001556020105774300007c3a00001582020105ba0300000941000015bb03010591060000f50d000015120601001d68800100000000000e0000000152023f000058390000158b0703111a1900006a800100000000000c000000158c0705090e1900006a800100000000000c000000048605000000026948000002ff430000058d2d0000b94600001be40401058d2d0000b94600001be404010529460000594b00001bcd04010529460000594b00001bcd0401000002cb190000023c260000153680010000000000120000000152bf440000933000001ebb0211721000003680010000000000120000001ebc021b11371300003680010000000000120000000944070909651000003680010000000000120000001f591200000000021c320000154880010000000000120000000152c2020000933000001ed60211721000004880010000000000120000001ed7021b11371300004880010000000000120000000944070909651000004880010000000000120000001f5912000000000002fb130000035a800100000000000e0000000152ec0400001e12000020720602714700000531320000a71800002025050105cd060000d73b00002025050100024130000005923e00005b090000209b07010000029126000002e7170000058a220000b02b000022580101058a220000b02b0000225801010002413000000e6486010000000000a200000001522e1000009330000022830f62110000f00c000022830a12f9160000200d000009e6071b0c65100000500d00001f1701120011c1160000a2860100000000005800000009e807091168210000ac860100000000004a0000001f65012711b5150000ae86010000000000480000002027051611c9150000c286010000000000060000001f66013c0bc9040000c286010000000000060000001f700109000b65100000ca86010000000000140000001f6701150b65100000e086010000000000160000001f69011100000000000000028c060000020335000005022d000030180000269906010539180000352d000026b50601029730000005731500007c4400002677020100000000002c0000000200000000000800ffffffffe8420100000000000e0000000000000000000000000000000000000000000000bc0100000200510000000800ffffffffa2770100000000000400000000000000a6770100000000000e00000000000000b4770100000000000200000000000000b6770100000000004201000000000000f878010000000000e401000000000000dc7a0100000000005600000000000000327b0100000000007803000000000000aa7e0100000000000e00000000000000b87e0100000000007e0100000000000036800100000000001200000000000000488001000000000012000000000000005a800100000000000e0000000000000068800100000000000e0000000000000076800100000000007000000000000000e680010000000000bc01000000000000a282010000000000b400000000000000568301000000000038000000000000008e830100000000000a000000000000009883010000000000b6000000000000004e840100000000003a0000000000000088840100000000002001000000000000a885010000000000980000000000000040860100000000000e000000000000004e8601000000000016000000000000006486010000000000a200000000000000068701000000000070000000000000000000000000000000000000000000000028780100000000002c780100000000003078010000000000387801000000000044780100000000004878010000000000000000000000000000000000000000003a780100000000004278010000000000487801000000000050780100000000000000000000000000000000000000000082780100000000008e7801000000000090780100000000009a7801000000000000000000000000000000000000000000bc78010000000000c878010000000000ca78010000000000d27801000000000000000000000000000000000000000000727901000000000078790100000000007c790100000000008279010000000000367a010000000000667a01000000000000000000000000000000000000000000967a010000000000b67a010000000000d67a010000000000dc7a010000000000000000000000000000000000000000009e7a010000000000a67a010000000000d67a010000000000dc7a010000000000000000000000000000000000000000009e7a010000000000a67a010000000000d67a010000000000dc7a010000000000000000000000000000000000000000009e7a010000000000a67a010000000000d67a010000000000dc7a01000000000000000000000000000000000000000000e879010000000000ee79010000000000fc79010000000000007a01000000000000000000000000000000000000000000ee79010000000000f279010000000000007a010000000000047a0100000000000000000000000000000000000000000044790100000000004879010000000000507901000000000052790100000000005a790100000000005c790100000000005e7901000000000060790100000000000000000000000000000000000000000052790100000000005a790100000000005c790100000000005e7901000000000000000000000000000000000000000000347b0100000000004a7b0100000000004c7b010000000000547b01000000000000000000000000000000000000000000347b0100000000004a7b0100000000004c7b010000000000547b01000000000000000000000000000000000000000000767b010000000000807b010000000000887b010000000000d27b01000000000000000000000000000000000000000000767b0100000000007a7b010000000000887b010000000000ce7b01000000000000000000000000000000000000000000767b0100000000007a7b010000000000887b010000000000ce7b010000000000000000000000000000000000000000003e7c010000000000547c0100000000005a7c0100000000005e7c010000000000000000000000000000000000000000003e7c010000000000547c0100000000005a7c0100000000005e7c01000000000000000000000000000000000000000000567c0100000000005a7c010000000000607c010000000000627c01000000000000000000000000000000000000000000787c0100000000007c7c010000000000847c010000000000867c0100000000008e7c010000000000907c010000000000927c010000000000967c01000000000000000000000000000000000000000000867c0100000000008e7c010000000000907c010000000000927c01000000000000000000000000000000000000000000aa7c010000000000ae7c010000000000b47c010000000000b67c010000000000be7c010000000000c07c010000000000c27c010000000000c47c01000000000000000000000000000000000000000000b67c010000000000be7c010000000000c07c010000000000c27c01000000000000000000000000000000000000000000c67c010000000000c87c010000000000d27c010000000000d47c010000000000dc7c010000000000de7c010000000000e07c010000000000e27c01000000000000000000000000000000000000000000d47c010000000000dc7c010000000000de7c010000000000e07c010000000000000000000000000000000000000000004c7d0100000000004e7d010000000000927d010000000000967d010000000000987d0100000000009e7d01000000000000000000000000000000000000000000567d0100000000005e7d010000000000607d010000000000647d010000000000667d0100000000006c7d0100000000006e7d0100000000007e7d010000000000807d010000000000827d010000000000867d010000000000927d010000000000000000000000000000000000000000009e7d010000000000b67d010000000000b87d010000000000ba7d010000000000c67d010000000000c87d010000000000ca7d010000000000ce7d01000000000000000000000000000000000000000000e87d010000000000ee7d010000000000f27d010000000000f87d0100000000001e7e010000000000507e01000000000000000000000000000000000000000000747e0100000000007c7e0100000000008e7e010000000000927e01000000000000000000000000000000000000000000747e0100000000007c7e0100000000008e7e010000000000927e01000000000000000000000000000000000000000000747e010000000000787e0100000000008e7e010000000000927e01000000000000000000000000000000000000000000d07e010000000000d87e010000000000dc7e010000000000e47e01000000000000000000000000000000000000000000ea7e010000000000147f010000000000947f010000000000a47f01000000000000000000000000000000000000000000ea7e010000000000147f010000000000947f010000000000a47f01000000000000000000000000000000000000000000267f010000000000347f010000000000387f010000000000927f01000000000000000000000000000000000000000000a87f010000000000c67f010000000000e47f010000000000ee7f01000000000000000000000000000000000000000000a87f010000000000c67f010000000000e47f010000000000ee7f01000000000000000000000000000000000000000000f27f010000000000f87f010000000000fe7f010000000000028001000000000006800100000000000a8001000000000000000000000000000000000000000000f27f010000000000f87f010000000000fe7f010000000000028001000000000006800100000000000a80010000000000000000000000000000000000000000007c80010000000000d280010000000000d880010000000000e680010000000000000000000000000000000000000000008c800100000000008e80010000000000a480010000000000a88001000000000000000000000000000000000000000000b280010000000000bc80010000000000d880010000000000e68001000000000000000000000000000000000000000000b280010000000000bc80010000000000d880010000000000e68001000000000000000000000000000000000000000000b280010000000000bc80010000000000d880010000000000e680010000000000000000000000000000000000000000002c81010000000000448101000000000064810100000000004082010000000000000000000000000000000000000000002c8101000000000044810100000000006481010000000000408201000000000000000000000000000000000000000000448101000000000052810100000000007082010000000000748201000000000000000000000000000000000000000000448101000000000052810100000000007082010000000000748201000000000000000000000000000000000000000000448101000000000052810100000000007082010000000000748201000000000000000000000000000000000000000000448101000000000052810100000000007082010000000000748201000000000000000000000000000000000000000000b082010000000000b482010000000000bc82010000000000c282010000000000de82010000000000e48201000000000000000000000000000000000000000000a883010000000000ac83010000000000b483010000000000ba83010000000000d683010000000000dc83010000000000000000000000000000000000000000009e84010000000000a084010000000000ac840100000000008a8501000000000000000000000000000000000000000000b084010000000000b484010000000000b884010000000000bc8401000000000000000000000000000000000000000000b084010000000000b484010000000000b884010000000000bc8401000000000000000000000000000000000000000000fa84010000000000048501000000000006850100000000000a850100000000000000000000000000000000000000000018850100000000001c850100000000002285010000000000608501000000000064850100000000006e850100000000000000000000000000000000000000000018850100000000001c850100000000002285010000000000608501000000000064850100000000006e85010000000000000000000000000000000000000000006e8601000000000070860100000000007286010000000000fa86010000000000000000000000000000000000000000006e86010000000000708601000000000072860100000000008e86010000000000000000000000000000000000000000006e86010000000000708601000000000072860100000000008286010000000000000000000000000000000000000000000c87010000000000628701000000000068870100000000007687010000000000000000000000000000000000000000001c870100000000001e87010000000000348701000000000038870100000000000000000000000000000000000000000042870100000000004c87010000000000688701000000000076870100000000000000000000000000000000000000000042870100000000004c87010000000000688701000000000076870100000000000000000000000000000000000000000042870100000000004c870100000000006887010000000000768701000000000000000000000000000000000000000000a277010000000000a677010000000000a677010000000000b477010000000000b477010000000000b677010000000000b677010000000000f878010000000000f878010000000000dc7a010000000000dc7a010000000000327b010000000000327b010000000000aa7e010000000000aa7e010000000000b87e010000000000b87e01000000000036800100000000003680010000000000488001000000000048800100000000005a800100000000005a800100000000006880010000000000688001000000000076800100000000007680010000000000e680010000000000e680010000000000a282010000000000a282010000000000568301000000000056830100000000008e830100000000008e83010000000000988301000000000098830100000000004e840100000000004e8401000000000088840100000000008884010000000000a885010000000000a885010000000000408601000000000040860100000000004e860100000000004e8601000000000064860100000000006486010000000000068701000000000006870100000000007687010000000000000000000000000000000000000000007261775f7665630073747200636f756e74005f5a4e34636f726535736c6963653469746572313349746572244c542454244754243134706f73745f696e635f73746172743137683231633736663939343638653065646545007b636c6f7375726523307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e005f5a4e34636f726533707472347265616431376831626239643039646638396234373532450077726974653c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e007b696d706c2335347d00616476616e63655f62793c636f72653a3a7374723a3a697465723a3a43686172496e64696365733e006e657874005f5a4e34636f726533737472367472616974733131305f244c5424696d706c2475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c5424737472244754242475323024666f722475323024636f72652e2e6f70732e2e72616e67652e2e52616e6765546f244c54247573697a652447542424475424336765743137683633326532303137643665353735396645006e6578743c5b7573697a653b20345d3e00636f6e7461696e735f6e6f6e5f636f6e74696e756174696f6e5f62797465006275696c64657273005f5a4e3131305f244c5424636f72652e2e6f70732e2e72616e67652e2e52616e676546726f6d244c54247573697a6524475424247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c54242475356224542475356424244754242447542435696e6465783137686163396536316662616530626263376145005f5a4e34636f726533666d7439466f726d617474657231327061645f696e74656772616c3137686238656639343965396131613633346545005f5a4e36335f244c5424636f72652e2e63656c6c2e2e426f72726f774d75744572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683636336332373865383138373636393045005f5a4e34636f726533666d74336e756d35335f244c5424696d706c2475323024636f72652e2e666d742e2e55707065724865782475323024666f7224753230246936342447542433666d743137683464336136353331313038303933376445005f5a4e34636f726533666d7439466f726d617474657239616c7465726e617465313768333537326537646636323036356664374500696e646578005f5a4e34636f7265366f7074696f6e31354f7074696f6e244c5424542447542439756e777261705f6f72313768343165333439646137383638346138334500616c69676e5f6f66667365743c75383e005f5a4e34636f72653373747232315f244c5424696d706c24753230247374722447542439656e64735f776974683137683139626662313333653233336465306145005f5a4e34636f726535736c69636532395f244c5424696d706c2475323024247535622454247535642424475424336765743137683233646638653962656438656665346645005f5a4e34636f726533666d74386275696c64657273313044656275675475706c65356669656c6432385f24753762242475376224636c6f73757265247537642424753764243137686363643963626231656235626135633645005f5a4e34636f726536726573756c743133756e777261705f6661696c65643137683030653934303161326339653536633045007074720070616464696e670077726974653c636861723e0069735f736f6d653c7573697a653e00676574005f5a4e37355f244c54247573697a65247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c542424753562245424753564242447542424475424336765743137683362336666656535366439303731313345005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243873706c69745f61743137683461343239666364306233623563343945005f5a4e3131305f244c5424636f72652e2e697465722e2e61646170746572732e2e656e756d65726174652e2e456e756d6572617465244c54244924475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e65787431376831623734616564656639323065303665450063686172005f5a4e34636f7265366f7074696f6e31354f7074696f6e244c5424542447542436696e736572743137686265366237313331636461646331646245005f5a4e34636f726536726573756c743139526573756c74244c542454244324452447542438616e645f7468656e313768316532623263316238653933626561654500636f70795f66726f6d5f736c696365005f5a4e34636f726533666d7439466f726d6174746572323564656275675f7475706c655f6669656c64315f66696e6973683137683963326264643732306464613133376545007b696d706c2332397d007b696d706c2336357d005f5a4e3130385f244c5424636f72652e2e697465722e2e61646170746572732e2e66696c7465722e2e46696c746572244c5424492443245024475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722447542435636f756e743137683631323362313132363938303130326445005f5a4e34636f72653370747235777269746531376830336462313664353065636536366165450072616e6765006f7074696f6e005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f72336e74683137683635613666633036633265613031396645005f5a4e34636f72653373747235636f756e743134646f5f636f756e745f6368617273313768653066306166323562653730356463664500616c69676e5f746f5f6f6666736574733c75382c207573697a653e005f5a4e34636f726533636d70336d696e3137683961303232643031326665326338333745007b696d706c23317d005f5a4e34636f726533666d743372756e313768666639613633333362396633663061614500676574636f756e7400697465725f6d75743c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e006272616e63683c28292c20636f72653a3a666d743a3a4572726f723e007b696d706c2332357d005f5a4e34636f7265336f70733866756e6374696f6e36466e4f6e63653963616c6c5f6f6e63653137683331326365396462383432326365623645005f5a4e34636f726533666d74386275696c64657273313044656275675475706c65356669656c643137686134393061356537663734366534656245005f5a4e34636f72653130696e7472696e736963733139636f70795f6e6f6e6f7665726c617070696e673137683165326664363834393232323263326345005f5a4e34636f726533666d7439466f726d6174746572397369676e5f706c75733137683765363563323535316433616561343445007369676e5f706c7573005f5a4e34636f72653373747235636f756e743233636861725f636f756e745f67656e6572616c5f6361736531376864313333363866323830386530613030450076616c69646174696f6e73005f5a4e34636f726535736c696365346974657238375f244c5424696d706c2475323024636f72652e2e697465722e2e7472616974732e2e636f6c6c6563742e2e496e746f4974657261746f722475323024666f7224753230242452462424753562245424753564242447542439696e746f5f697465723137683765326332623733366531386264656545005f5a4e34636f726533707472376d75745f70747233315f244c5424696d706c2475323024244250246d75742475323024542447542433616464313768333939313037663564323335643062374500497465724d75740047656e657269635261646978006e6578745f696e636c75736976653c636861723e005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243132616c69676e5f6f66667365743137686265366661383332613635626436303545007b696d706c2335337d0064726f705f696e5f706c6163653c26636f72653a3a697465723a3a61646170746572733a3a636f706965643a3a436f706965643c636f72653a3a736c6963653a3a697465723a3a497465723c75383e3e3e005f5a4e34636f7265337074723133726561645f766f6c6174696c653137683034656338646164326362346562306245006d75745f7074720073756d005f5a4e34636f726533666d7439466f726d61747465723770616464696e67313768386664646163386139653836623737364500636d7000696d706c73005f5a4e34636f72653373747232315f244c5424696d706c247532302473747224475424313669735f636861725f626f756e646172793137683034353265303532643135616334353245005f5a4e37355f244c54247573697a65247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c542424753562245424753564242447542424475424336765743137686337356165633633323166633531643545005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542439656e64735f77697468313768383363653331633938643238356662364500696e736572743c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e005f5a4e34636f72653970616e69636b696e673970616e69635f666d743137686436616161656662346334646538633945005f5a4e34636f72653373747235636f756e743131636f756e745f63686172733137683362393037393633646461313835376345007265706c6163653c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e005f5a4e34636f7265366f7074696f6e31354f7074696f6e244c542454244754243769735f736f6d653137686166353061376333383437653666373645006e74683c636f72653a3a7374723a3a697465723a3a43686172496e64696365733e005f5a4e34636f726533737472313176616c69646174696f6e733135757466385f66697273745f627974653137683962396637633933306431356335663945005f5a4e34636f726533666d7438676574636f756e743137683639663830313763343363306364653245005f5a4e34636f72653970616e69636b696e673970616e69635f7374723137683666303932373830653338346562353045005f5a4e34636f726535736c696365366d656d6368723138636f6e7461696e735f7a65726f5f627974653137686130353638656531383330306135373245005f5a4e34355f244c5424244c502424525024247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d74313768613430323766643039663261636331324500666d743c28293e005f5a4e36375f244c5424636f72652e2e61727261792e2e54727946726f6d536c6963654572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d74313768353264643636336235383463633535664500636f70795f6e6f6e6f7665726c617070696e673c75383e00616363756d007b696d706c2334387d007b636c6f7375726523307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542434697465723137686266616536663139613561623764656445006765745f756e636865636b65643c636f72653a3a666d743a3a72743a3a417267756d656e742c207573697a653e006765743c267374723e0070616e69635f646973706c61793c267374723e00756e777261705f6661696c6564002f72757374632f32663662633564323539653761623235646466646433336465353362383932373730323138393138007274005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f7234666f6c64313768623061333862663336373733633236364500636f756e743c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e005f5a4e34636f726533707472347265616431376831653634383335653639376533366630450073756d5f62797465735f696e5f7573697a65005f5a4e34636f726533666d7432727438417267756d656e743861735f7573697a653137686437613231613332353662616362386245005f5a4e3131305f244c5424636f72652e2e697465722e2e61646170746572732e2e656e756d65726174652e2e456e756d6572617465244c54244924475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e657874313768633030313137313163643937383139624500726573756c74005f5a4e37335f244c5424636f72652e2e666d742e2e6e756d2e2e4c6f776572486578247532302461732475323024636f72652e2e666d742e2e6e756d2e2e47656e657269635261646978244754243564696769743137686634306237613733623764393162653445004d61796265556e696e6974007b696d706c2336347d005f5a4e37335f244c54242475356224412475356424247532302461732475323024636f72652e2e736c6963652e2e636d702e2e536c6963655061727469616c4571244c542442244754242447542435657175616c3137686637383434376536346661643333376145005f5a4e3130365f244c5424636f72652e2e6f70732e2e72616e67652e2e52616e6765244c54247573697a6524475424247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c542424753562245424753564242447542424475424336765743137683761383664333261616263343034303345005f5a4e34636f72653463686172376d6574686f647332325f244c5424696d706c247532302463686172244754243131656e636f64655f757466383137683661333732316366346263313738623645005f5a4e34636f726533666d74336e756d33696d7037666d745f7536343137683238366534643532373433386334363745005f5a4e34636f72653970616e69636b696e673570616e69633137686437373538656430613265383739363145006c6962726172792f636f72652f7372632f6c69622e72732f402f636f72652e353431663036343835316338633866372d6367752e3000726561645f766f6c6174696c653c7573697a653e005f5a4e3130385f244c5424636f72652e2e697465722e2e61646170746572732e2e66696c7465722e2e46696c746572244c5424492443245024475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722447542435636f756e7438746f5f7573697a6532385f24753762242475376224636c6f73757265247537642424753764243137686532646263323632336436376436643345005f5a4e34636f726533666d743131506f737450616464696e673577726974653137683130373832303864313037663934393045006164643c7573697a653e005f5a4e34636f726533666d7439466f726d61747465723977726974655f737472313768353330393765363135313339346565644500696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e2c20636f72653a3a6f70733a3a72616e67653a3a52616e676546726f6d3c7573697a653e3e007b696d706c2331357d00656e64735f776974683c75383e005f5a4e34636f726535736c696365366d656d636872366d656d6368723137683838333063653264646237323666636245006c656e5f75746638005f5a4e34636f72653463686172376d6574686f64733135656e636f64655f757466385f7261773137686230336466376165346464366562316445005f5a4e34636f726533666d74355772697465313077726974655f63686172313768666466623438666364333637346132384500616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23347d3a3a6669656c643a3a7b636c6f737572655f656e7623307d3e00636f7265005f5a4e34636f726533636d7035696d706c7335375f244c5424696d706c2475323024636f72652e2e636d702e2e5061727469616c4f72642475323024666f7224753230247573697a6524475424326c74313768383563303932356636663163316566654500646f5f636f756e745f6368617273005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542431336765745f756e636865636b656431376838333832313033623533356331333034450063656c6c006765743c75382c20636f72653a3a6f70733a3a72616e67653a3a52616e67653c7573697a653e3e0066696e6973680077726974655f70726566697800636861725f636f756e745f67656e6572616c5f6361736500706f73745f696e635f73746172743c75383e007265706c6163653c636861723e00506f737450616464696e6700697465723c75383e005f5a4e38375f244c5424636f72652e2e7374722e2e697465722e2e43686172496e6469636573247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683862646365633661316137393933386345005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542433676574313768396431656137353833353464396166364500656e756d6572617465005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683563636236663439653430616432356245005f5a4e34636f726535736c69636534697465723136497465724d7574244c54245424475424336e65773137683131393134666634646337396132326545006469676974005f5a4e34636f726535736c69636533636d7038315f244c5424696d706c2475323024636f72652e2e636d702e2e5061727469616c4571244c54242475356224422475356424244754242475323024666f7224753230242475356224412475356424244754243265713137683331383339323064643563373930336445006d656d6368725f616c69676e656400777261705f6275663c636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23317d3a3a777261703a3a7b636c6f737572655f656e7623307d3e005f5a4e34636f726533666d74386275696c6465727331305061644164617074657234777261703137686630613261643433323636313138356545005f5a4e34636f726533666d74386275696c64657273313044656275675475706c653666696e6973683137683262326465366164386361323965353845006974657200666f6c643c7573697a652c20636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c207573697a652c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e005f5a4e34636f72653373747235636f756e743233636861725f636f756e745f67656e6572616c5f6361736532385f24753762242475376224636c6f73757265247537642424753764243137686238333838383631636166343538396545007b636c6f7375726523307d3c2675382c207573697a652c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e00737065635f6e6578743c7573697a653e005f5a4e34636f726534697465723572616e67653130315f244c5424696d706c2475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722475323024666f722475323024636f72652e2e6f70732e2e72616e67652e2e52616e6765244c5424412447542424475424346e6578743137683166316635393732633862353338396245005f5a4e34636f726533737472313176616c69646174696f6e733138757466385f6163635f636f6e745f62797465313768386431353839303565613233346333334500757466385f6163635f636f6e745f62797465006164643c5b7573697a653b20345d3e006e65773c5b7573697a653b20345d3e005f5a4e34636f726535736c6963653469746572313349746572244c542454244754243134706f73745f696e635f73746172743137686632323465323937613136633263656145006e6578743c636f72653a3a736c6963653a3a697465723a3a497465723c636f72653a3a666d743a3a72743a3a417267756d656e743e3e005f5a4e34636f726535617272617938355f244c5424696d706c2475323024636f72652e2e6f70732e2e696e6465782e2e496e646578244c542449244754242475323024666f722475323024247535622454247533622424753230244e24753564242447542435696e6465783137683663646534633833393961376530333445007b696d706c23397d0064656275675f7475706c655f6e6577005f5a4e34636f726533666d74386275696c64657273313044656275675475706c653666696e69736832385f24753762242475376224636c6f737572652475376424247537642431376861393666623161373161643166373535450064656275675f7475706c655f6669656c64315f66696e697368006164643c75383e007b696d706c233138317d00666f6c643c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a6d61703a3a6d61705f666f6c643a3a7b636c6f737572655f656e7623307d3c2675382c207573697a652c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e3e005f5a4e34636f726535736c69636532395f244c5424696d706c2475323024247535622454247535642424475424313873706c69745f61745f756e636865636b65643137683765396534313435376636393734393145006e6578743c636f72653a3a736c6963653a3a697465723a3a497465723c636f72653a3a666d743a3a72743a3a506c616365686f6c6465723e3e007b696d706c2331377d005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542438697465725f6d75743137683030376635633136366631613761373245006172726179005f5a4e34636f7265337374723469746572323253706c6974496e7465726e616c244c5424502447542431346e6578745f696e636c75736976653137683938613230353930343932666138366445005f5a4e35325f244c542463686172247532302461732475323024636f72652e2e7374722e2e7061747465726e2e2e5061747465726e24475424313269735f7375666669785f6f663137683866653837336364343736333664316445005f5a4e34636f726533666d7439466f726d617474657238777261705f6275663137686636336162363038633262616362303045007b636c6f7375726523307d0070616e69636b696e67005f5a4e35365f244c54247573697a65247532302461732475323024636f72652e2e697465722e2e7472616974732e2e616363756d2e2e53756d244754243373756d3137683739356164323965353439386433333445005f5a4e34636f72653373747232315f244c5424696d706c2475323024737472244754243132636861725f696e64696365733137686466343535663065643137623532303045006765743c75382c207573697a653e005f5a4e34636f7265337074723132616c69676e5f6f66667365743137683534623332333739346162326331313545005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243961735f6368756e6b7331376831643562356538303063366463326238450061735f6368756e6b733c7573697a652c20343e005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e737424753230245424475424336164643137683566666465653639383065666566633145006765745f756e636865636b65643c636f72653a3a666d743a3a72743a3a417267756d656e743e0064656275675f737472756374007b696d706c2332387d0065713c5b75385d2c205b75385d3e0044656275675475706c6500666d745f696e743c636f72653a3a666d743a3a6e756d3a3a55707065724865782c207536343e00636c616e67204c4c564d202872757374632076657273696f6e20312e37312e302d6e696768746c79202832663662633564323520323032332d30352d30392929006974657261746f72005f5a4e34636f726533737472313176616c69646174696f6e7331356e6578745f636f64655f706f696e74313768656364656330303032323838613566354500757466385f66697273745f627974650069735f636861725f626f756e64617279006d696e3c7573697a653e005f5a4e34636f72653373747235636f756e743330636f6e7461696e735f6e6f6e5f636f6e74696e756174696f6e5f627974653137686530636638653465356130663030393045005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137686134633765313364663063343439373145005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243361646431376833356564316564666234363437623138450077726974655f737472005f5a4e34636f726533666d74336e756d313247656e65726963526164697837666d745f696e743137686162643431393537653230363731373445006d617962655f756e696e697400696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e2c20636f72653a3a6f70733a3a72616e67653a3a52616e676546726f6d3c7573697a653e2c203132383e005f5a4e39395f244c5424636f72652e2e7374722e2e697465722e2e53706c6974496e636c7573697665244c54245024475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683536356238663563313134366339666645005f5a4e38315f244c5424636f72652e2e7374722e2e7061747465726e2e2e436861725365617263686572247532302461732475323024636f72652e2e7374722e2e7061747465726e2e2e53656172636865722447542431306e6578745f6d617463683137686231353436643361613035653433333145005f5a4e34636f72653463686172376d6574686f6473386c656e5f75746638313768343935363635353564666635366333654500656e636f64655f757466385f72617700616c6c6f6300747261697473005f5a4e34636f726535736c6963653469746572313349746572244c54245424475424336e65773137683436326338393130346236666239373745005f5a4e34636f7265336e756d32335f244c5424696d706c24753230247573697a652447542431327772617070696e675f6d756c3137683933396664623563663661656266303945006e6577006d656d6368720077726170005f5a4e34636f726533666d74336e756d313247656e65726963526164697837666d745f696e743137683330323730653937613764383866626145007061640070616e6963005f5a4e34636f726533666d74336e756d35335f244c5424696d706c2475323024636f72652e2e666d742e2e4c6f7765724865782475323024666f7224753230246936342447542433666d74313768663235653065383534373535336437314500696d7000616c7465726e617465006d6170005f5a4e3130325f244c5424636f72652e2e697465722e2e61646170746572732e2e6d61702e2e4d6170244c5424492443244624475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722447542434666f6c643137683439653563633739303661396231626645007772697465007b696d706c23377d006d696e5f62793c7573697a652c20666e28267573697a652c20267573697a6529202d3e20636f72653a3a636d703a3a4f72646572696e673e006765743c267374722c207573697a653e005f5a4e34636f726535736c69636535696e64657837345f244c5424696d706c2475323024636f72652e2e6f70732e2e696e6465782e2e496e646578244c542449244754242475323024666f72247532302424753562245424753564242447542435696e64657831376835623336343435386238326632343635450053706c6974496e7465726e616c006e6578743c636861723e0057726974650077726974655f636861723c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e007b696d706c2332367d005f5a4e34325f244c54242452462454247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d74313768633230363132656137383639386165344500666d74007b696d706c23307d004f7074696f6e007b696d706c23387d005f5a4e34636f726533707472376d75745f70747233315f244c5424696d706c2475323024244250246d757424753230245424475424336164643137686433383935323761353331303836366545006765745f756e636865636b65643c267374723e005f5a4e34636f726533666d7439466f726d6174746572313264656275675f73747275637431376838333134343030643138313466376534450070616e69635f737472005f5a4e34636f726533666d74386275696c64657273313564656275675f7475706c655f6e65773137683134383664383033383865636636373745005553495a455f4d41524b455200736c696365005f5a4e34636f7265336d656d377265706c6163653137683665313530623565366261663964346545007061645f696e74656772616c006765743c75383e005f5a4e34636f726535736c6963653469746572313349746572244c54245424475424336e65773137686231373834333338323430613463363745007b696d706c2331397d006e6578745f6d61746368005f5a4e34636f726536726573756c743139526573756c74244c542454244324452447542438616e645f7468656e3137686639613762303833656534636237383245005f5a4e37335f244c5424636f72652e2e666d742e2e6e756d2e2e5570706572486578247532302461732475323024636f72652e2e666d742e2e6e756d2e2e47656e657269635261646978244754243564696769743137683933663339316566393536306361643245005f5a4e34636f72653370747231303264726f705f696e5f706c616365244c542424524624636f72652e2e697465722e2e61646170746572732e2e636f706965642e2e436f70696564244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c542475382447542424475424244754243137683465633534623435323134663763393045005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683334323336653433336537396333623345006c74006368617273005f5a4e34636f72653373747232315f244c5424696d706c247532302473747224475424336765743137686361316261643162613538333362626645006765743c636f72653a3a6f70733a3a72616e67653a3a52616e6765546f3c7573697a653e3e00706f73745f696e635f73746172743c7573697a653e005f5a4e37355f244c54247573697a65247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c54242475356224542475356424244754242447542431336765745f756e636865636b65643137686630663432666234656339376261626145006164643c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e006d6574686f6473005f5a4e34636f726533666d74386275696c64657273313050616441646170746572347772617032385f24753762242475376224636c6f737572652475376424247537642431376862353032353031383864353564626337450063617061636974795f6f766572666c6f7700666d745f753634005f5a4e36385f244c5424636f72652e2e666d742e2e6275696c646572732e2e50616441646170746572247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f7374723137686539366438303337316562386433343445005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243361646431376836343831303738333031643161616237450049746572005f5a4e34636f72653373747232315f244c5424696d706c2475323024737472244754243563686172733137683635643537336338666664393434333645005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f723130616476616e63655f62793137683837343136383366376333383664636245006e6578745f636f64655f706f696e743c636f72653a3a736c6963653a3a697465723a3a497465723c75383e3e005f5a4e39335f244c5424636f72652e2e736c6963652e2e697465722e2e4368756e6b73244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137686264343939663734373230663065386245004f7264006164643c267374723e007b696d706c23367d005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f666d743137683565373464633863623261616161323645007b696d706c23327d005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542434697465723137686331616261316236653465646465623545005f5a4e34636f726533666d7439466f726d6174746572336e65773137686165623034366666366431666231663445005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243361646431376838353436653232346135313966363633450064656275675f7374727563745f6e657700746f5f7538005f5a4e34636f726533636d7035696d706c7336395f244c5424696d706c2475323024636f72652e2e636d702e2e5061727469616c4571244c54242452462442244754242475323024666f7224753230242452462441244754243265713137683436393566636435376362636161326145005f5a4e34636f726533666d743577726974653137683537653362636463656237646630393145006578706563745f6661696c6564006c656e5f6d69736d617463685f6661696c006f707300696e7472696e736963730073756d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e005f5a4e34636f7265336d656d377265706c61636531376838363534306363336630326138396663450069735f6e6f6e653c7573697a653e00697465723c5b7573697a653b20345d3e00696e746f5f697465723c5b7573697a653b20345d3e005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683366313636623661373436326234373945005f5a4e34636f726533666d7432727438417267756d656e7433666d74313768363232636537653835383430326338654500666d745f696e743c636f72653a3a666d743a3a6e756d3a3a4c6f7765724865782c207536343e00657175616c3c75382c2075383e005f5a4e34636f726535736c696365366d656d63687231326d656d6368725f6e616976653137686363623962373463393862393633336245006d656d6368725f6e6169766500616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23347d3a3a66696e6973683a3a7b636c6f737572655f656e7623307d3e00636f6e73745f707472005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f723373756d313768616537613566613764646461346162384500757466385f69735f636f6e745f62797465006e6578743c636f72653a3a666d743a3a72743a3a417267756d656e743e005f5a4e34636f726533666d74386275696c64657273313664656275675f7374727563745f6e65773137686135363836656238343531653037323245005f5a4e34636f72653970616e69636b696e67313370616e69635f646973706c6179313768663965353336303933393038663832624500656e64735f776974683c636861723e0065713c75382c2075383e007b696d706c23347d005f5a4e34636f726533737472313176616c69646174696f6e733137757466385f69735f636f6e745f6279746531376861396331376363326537313134623836450073706c69745f61745f756e636865636b65643c75383e0073706c69745f61743c75383e005f5a4e34636f72653373747235636f756e74313873756d5f62797465735f696e5f7573697a653137683733663965326535343130353136333245006e6578743c636f72653a3a666d743a3a72743a3a506c616365686f6c6465723e00417267756d656e74005f5a4e37355f244c54247573697a65247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c54242475356224542475356424244754242447542431336765745f756e636865636b6564313768656630633435353430343632353962624500636f6e7461696e735f7a65726f5f62797465005f5a4e37395f244c5424636f72652e2e726573756c742e2e526573756c74244c5424542443244524475424247532302461732475323024636f72652e2e6f70732e2e7472795f74726169742e2e54727924475424366272616e63683137683034646133323232663535363066313845005f5a4e34636f7265366f7074696f6e31336578706563745f6661696c65643137686332333330616533386638616564396545005f5a4e34636f726533707472376d75745f70747233315f244c5424696d706c2475323024244250246d7574247532302454244754243361646431376837336363316163653933303039363536450073756d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e2c207573697a653e005f5a4e35365f244c54247573697a65247532302461732475323024636f72652e2e697465722e2e7472616974732e2e616363756d2e2e53756d244754243373756d32385f24753762242475376224636c6f73757265247537642424753764243137683665653564323561643365666465373945007369676e5f61776172655f7a65726f5f70616400726561643c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e006e6578743c7573697a653e00756e777261705f6f723c267374723e005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243136616c69676e5f746f5f6f6666736574733137683265333033653231353164623038353745005f5a4e34636f726535736c69636532395f244c5424696d706c2475323024247535622454247535642424475424336765743137683037666466393631613031323632356145006e65773c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e007b696d706c2334347d0077726974655f7374723c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e577269746524475424313077726974655f636861723137683239666437616639333939643762333645005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243135636f70795f66726f6d5f736c69636531376c656e5f6d69736d617463685f6661696c3137686531663934356265353831313135613845006c6962726172792f616c6c6f632f7372632f6c69622e72732f402f616c6c6f632e643733613839653266303538366464312d6367752e30004974657261746f7200636f756e745f6368617273005f5a4e34636f72653469746572386164617074657273336d6170386d61705f666f6c6432385f24753762242475376224636c6f73757265247537642424753764243137686265643362346664336632356561633645005f5a4e34636f7265366f7074696f6e31354f7074696f6e244c542454244754243769735f6e6f6e653137683036303537623832613939663564313445005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542438616c69676e5f746f3137686361663565313535373365303734303345007b696d706c2331317d005f5a4e34636f726533636d70366d696e5f62793137683961363365346463336265666132393045005f5a4e34636f7265336d656d31326d617962655f756e696e697432304d61796265556e696e6974244c54245424475424357772697465313768643262633963366561386361383161624500656e636f64655f75746638005f5a4e34636f726533666d743557726974653977726974655f666d743137683364623431343565346436363932376245006669656c64005f5a4e36305f244c5424636f72652e2e63656c6c2e2e426f72726f774572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137686163386261333334363731373261333845006e6578743c75383e00746f5f7573697a65006d656d005f5a4e34636f7265337074723577726974653137683934303032343231393363646338316545005f5a4e38395f244c5424636f72652e2e6f70732e2e72616e67652e2e52616e6765244c54245424475424247532302461732475323024636f72652e2e697465722e2e72616e67652e2e52616e67654974657261746f72496d706c2447542439737065635f6e65787431376834303038636235396134653064623339450061735f7573697a65006164643c636f72653a3a666d743a3a72743a3a417267756d656e743e00696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e005f5a4e34636f7265336e756d32335f244c5424696d706c24753230247573697a652447542431327772617070696e675f73756231376838643635306338643866353735643162450069735f70726574747900616461707465727300726561643c636861723e007b696d706c23337d00636861725f696e646963657300616c69676e5f746f3c75382c207573697a653e007772617070696e675f6d756c0077726974653c75383e005f5a4e35305f244c5424753634247532302461732475323024636f72652e2e666d742e2e6e756d2e2e446973706c6179496e742447542435746f5f75383137683636316463333963356464386666653545007061747465726e0069735f7375666669785f6f66005f5a4e34636f726535736c696365366d656d63687231346d656d6368725f616c69676e6564313768643864383232303663636532343531614500526573756c7400506164416461707465720070616e69635f666d74005f5a4e34636f726533666d7439466f726d6174746572337061643137683433336537613934646232626438653245005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f7374723137683865303931326361326264646233386345005f5a4e34636f726533666d7432727431325553495a455f4d41524b455232385f24753762242475376224636c6f7375726524753764242475376424313768643137376134333532613130653633314500466e4f6e6365006e756d005f5a4e38315f244c5424636f72652e2e7374722e2e697465722e2e4368617273247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722447542435636f756e743137686638633866336432633063356164333545005f5a4e34636f726533666d7439466f726d617474657231397369676e5f61776172655f7a65726f5f7061643137683136323439616566366630343733333545006e65773c75383e007b696d706c23357d005f5a4e34636f726533636d70334f7264336d696e31376861623865636338303366663033636364450072756e005f5a4e34636f726533666d74386275696c64657273313044656275675475706c653969735f7072657474793137683131646663373739346165376162303045005f5a4e34636f726533666d7439466f726d617474657231327061645f696e74656772616c313277726974655f70726566697831376838346635386564303837613362643933450066756e6374696f6e00466f726d61747465720066696c746572006d61705f666f6c64005f5a4e38315f244c5424636f72652e2e7374722e2e697465722e2e4368617273247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683064323235303663643135633337363345007b696d706c2337307d005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683634663237353939353136663335636545005f5a4e35355f244c542424524624737472247532302461732475323024636f72652e2e7374722e2e7061747465726e2e2e5061747465726e24475424313269735f7375666669785f6f663137686536396533336230613062663235373545007772617070696e675f7375620077726974655f666d743c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e005f5a4e35616c6c6f63377261775f766563313763617061636974795f6f766572666c6f7731376837363964333737343539393364316265450063616c6c5f6f6e63653c636f72653a3a666d743a3a72743a3a5553495a455f4d41524b45523a3a7b636c6f737572655f656e7623307d2c2028267573697a652c20266d757420636f72653a3a666d743a3a466f726d6174746572293e003a000000020000000000510000003400000063617061636974795f6f766572666c6f77002f0000007261775f766563002a000000616c6c6f630000000000d51a0000020051000000ca2200006a01000077726974653c636861723e00161f00006d617962655f756e696e6974007b2100006272616e63683c28292c20636f72653a3a666d743a3a4572726f723e00e90000006d75745f70747200da1f0000696e736572743c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e0053190000636f70795f6e6f6e6f7665726c617070696e673c75383e00b7040000466f726d617474657200742000007b696d706c2331377d00001d0000737065635f6e6578743c7573697a653e00d6190000706f73745f696e635f73746172743c7573697a653e00381800007b696d706c2332357d0056210000526573756c74001b1e00006e6578745f636f64655f706f696e743c636f72653a3a736c6963653a3a697465723a3a497465723c75383e3e0034000000726561645f766f6c6174696c653c7573697a653e007b1a0000697465723c5b7573697a653b20345d3e00091f00007265706c6163653c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e00c11c00007b636c6f7375726523307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e00471a000073706c69745f61745f756e636865636b65643c75383e00fc1e00007265706c6163653c636861723e00c01f000069735f6e6f6e653c7573697a653e00951a00006765743c267374722c207573697a653e00af2100007b696d706c2332367d00771e000069735f636861725f626f756e646172790037210000726573756c74008718000066756e6374696f6e00b71c0000636f756e7400f00400007061645f696e74656772616c00611a0000616c69676e5f746f5f6f6666736574733c75382c207573697a653e00db1a00006c656e5f6d69736d617463685f6661696c00da0000006164643c75383e00be1900006e65773c75383e00e203000064696769740050180000666d743c28293e00d718000070616e69636b696e6700cd1f0000756e777261705f6f723c267374723e00951d0000636f6e7461696e735f6e6f6e5f636f6e74696e756174696f6e5f6279746500cd000000616c69676e5f6f66667365743c75383e000d1a00006e65773c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e00d52000007b696d706c2331397d00602000007772617070696e675f73756200c9040000616c7465726e617465004c1f00006c74008e1c00006d61705f666f6c6400a11d000073756d5f62797465735f696e5f7573697a6500ae010000417267756d656e74001b1f00004d61796265556e696e697400f4030000666d7400e81f00006578706563745f6661696c656400ef1b0000636f6e7461696e735f7a65726f5f6279746500a911000072756e00f61d00007b696d706c2334347d00bc1e00007b696d706c2332387d008d11000077726974655f707265666978008c180000466e4f6e636500261b00006765743c267374723e005b000000636f6e73745f70747200e71e00006e6578745f6d6174636800c91a00006765743c75382c20636f72653a3a6f70733a3a72616e67653a3a52616e67653c7573697a653e3e002d1f000077726974653c75383e00340100006164643c7573697a653e00ad19000049746572003713000064656275675f7374727563745f6e6577004b1800007b696d706c2335337d00b30000006164643c636f72653a3a666d743a3a72743a3a417267756d656e743e003d1d0000737472000e19000070616e69635f646973706c61793c267374723e00201a0000697465723c75383e00d61a0000636f70795f66726f6d5f736c69636500771c00006d617000b71e00007061747465726e00d9020000666d745f696e743c636f72653a3a666d743a3a6e756d3a3a4c6f7765724865782c207536343e00b015000066696e69736800dd0300007b696d706c2332397d0068210000616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23347d3a3a66696e6973683a3a7b636c6f737572655f656e7623307d3e003c210000756e777261705f6661696c656400701900006e6578743c75383e00e31d000053706c6974496e7465726e616c00711d0000646f5f636f756e745f636861727300a01900006e6578743c636f72653a3a666d743a3a72743a3a417267756d656e743e0061190000736c69636500c415000044656275675475706c6500bc1c0000746f5f7573697a6500b2190000706f73745f696e635f73746172743c75383e00ae1d000069746572005d1c000073756d00471f00007b696d706c2335347d00e31900007b696d706c2337307d001a1b00006765745f756e636865636b65643c636f72653a3a666d743a3a72743a3a417267756d656e743e00841700007b696d706c23307d005f1d0000636861725f636f756e745f67656e6572616c5f6361736500d41e000069735f7375666669785f6f6600811c0000666f6c643c7573697a652c20636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c207573697a652c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e007f100000777261705f6275663c636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23317d3a3a777261703a3a7b636c6f737572655f656e7623307d3e000918000077726974655f666d743c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e00e3010000666d745f753634002a000000636f7265006e1a000061735f6368756e6b733c7573697a652c20343e006211000064656275675f7475706c655f6669656c64315f66696e697368009c0100005553495a455f4d41524b455200721c0000616461707465727300462000007772617070696e675f6d756c00621c00007b636c6f7375726523307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e00831e00006765743c636f72653a3a6f70733a3a72616e67653a3a52616e6765546f3c7573697a653e3e00a60000006164643c5b7573697a653b20345d3e00ab1c0000636f756e743c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e00fb190000696e746f5f697465723c5b7573697a653b20345d3e00111c0000666f6c643c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a6d61703a3a6d61705f666f6c643a3a7b636c6f737572655f656e7623307d3c2675382c207573697a652c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e3e00e11600007b696d706c23317d008f2200006368617200a11c000066696c74657200d11c0000656e756d657261746500cb1b00006d656d6368725f6e6169766500dc18000070616e69635f666d7400e304000070616464696e6700160300007b696d706c2336347d004c1c00007b696d706c2334387d00e61600007772617000f916000064656275675f7475706c655f6e657700431300007b696d706c23327d00b301000061735f7573697a6500511c000073756d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e00421f0000696d706c7300471c0000616363756d0007170000577269746500f518000070616e696300941900006e6578743c636f72653a3a666d743a3a72743a3a506c616365686f6c6465723e005d1e0000636861727300821800006f707300942200006d6574686f647300ac1b000065713c75382c2075383e00fb1d00006e6578743c636861723e00ef0300007b696d706c2336357d00901e0000656e64735f776974683c636861723e00f71e00006d656d00cf1e00007b696d706c23337d001a19000070616e69635f73747200d61500006669656c6400881f00004f72640097010000727400de010000696d7000db1c00006e6578743c636f72653a3a736c6963653a3a697465723a3a497465723c636f72653a3a666d743a3a72743a3a506c616365686f6c6465723e3e00881900006e6578743c7573697a653e00081a0000497465724d757400c3110000777269746500af1a0000656e64735f776974683c75383e00c915000069735f707265747479007c1900006e6578743c5b7573697a653b20345d3e00e5020000666d745f696e743c636f72653a3a666d743a3a6e756d3a3a55707065724865782c207536343e002b1c0000616476616e63655f62793c636f72653a3a7374723a3a697465723a3a43686172496e64696365733e00d402000047656e657269635261646978009e1e0000747261697473008917000077726974655f7374723c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e00d61d00006e657874001e1c000073756d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e2c207573697a653e00981500007b696d706c23347d004813000077726974655f73747200992200006c656e5f75746638006c1f000065713c5b75385d2c205b75385d3e005d010000726561643c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e00541a000073706c69745f61743c75383e00e81d00006e6578745f696e636c75736976653c636861723e00040300007b696d706c2331317d0050010000726561643c636861723e00d907000070616400931c00007b636c6f7375726523307d3c2675382c207573697a652c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e00a217000077726974655f636861723c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e00271e0000757466385f66697273745f6279746500891b00007b696d706c23357d00e71c00006e6578743c636f72653a3a736c6963653a3a697465723a3a497465723c636f72653a3a666d743a3a72743a3a417267756d656e743e3e007b1f00006d696e5f62793c7573697a652c20666e28267573697a652c20267573697a6529202d3e20636f72653a3a636d703a3a4f72646572696e673e00591000006e6577002f2000006e756d007701000077726974653c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e00041b0000696e64657800ae1f00004f7074696f6e00b31f000069735f736f6d653c7573697a653e00321300006275696c64657273006a1e0000636861725f696e6469636573006f20000063656c6c00c00000006164643c267374723e002d1a00006765743c75382c207573697a653e003f1b00007b696d706c23367d00751b00006765743c75383e00b51500007b636c6f7375726523307d000f1e0000757466385f69735f636f6e745f62797465000c1c00004974657261746f72009118000063616c6c5f6f6e63653c636f72653a3a666d743a3a72743a3a5553495a455f4d41524b45523a3a7b636c6f737572655f656e7623307d2c2028267573697a652c20266d757420636f72653a3a666d743a3a466f726d6174746572293e00d71b00006d656d6368725f616c69676e6564003a1a0000616c69676e5f746f3c75382c207573697a653e00881a00006765745f756e636865636b65643c636f72653a3a666d743a3a72743a3a417267756d656e742c207573697a653e00410100006164643c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e00f61a0000697465725f6d75743c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e00a91f00006f7074696f6e00a6220000656e636f64655f757466385f726177000a1e000076616c69646174696f6e7300841b0000636d7000a81e000067657400321b00006765745f756e636865636b65643c267374723e00831100007b696d706c23377d006b1900007b696d706c233138317d00071c00006974657261746f72007210000064656275675f73747275637400631b0000696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e2c20636f72653a3a6f70733a3a72616e67653a3a52616e676546726f6d3c7573697a653e3e00381c00006e74683c636f72653a3a7374723a3a697465723a3a43686172496e64696365733e00b8220000656e636f64655f7574663800cf1600005061644164617074657200bf1b00006d656d63687200a31e00007b696d706c23387d0027190000696e7472696e7369637300a1210000696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e2c20636f72653a3a6f70733a3a72616e67653a3a52616e676546726f6d3c7573697a653e2c203132383e00f61c000072616e6765008f2100007b696d706c2331357d00d60400007369676e5f61776172655f7a65726f5f70616400bc0400007369676e5f706c7573002f000000707472004100000064726f705f696e5f706c6163653c26636f72653a3a697465723a3a61646170746572733a3a636f706965643a3a436f706965643c636f72653a3a736c6963653a3a697465723a3a497465723c75383e3e3e00531d0000636f756e745f636861727300ca1900006e65773c5b7573697a653b20345d3e0070110000506f737450616464696e67004b1e0000757466385f6163635f636f6e745f6279746500441b0000696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e005a1f00007b696d706c23397d00b6110000676574636f756e74005b210000616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23347d3a3a6669656c643a3a7b636c6f737572655f656e7623307d3e009b1f00006d696e3c7573697a653e0009030000746f5f7538008e1b0000657175616c3c75382c2075383e008a210000617272617900000000000e00000002000000000051000000000000000e000000020051000000ca22000000000000412a000000726973637600012000000004100572763634693270305f6d3270305f613270305f633270300058000000040034000000010101fb0e0d0001010101000000010000016c6962726172792f616c6c6f632f73726300007261775f7665632e72730001000000000902e842010000000000038a040105050a030109020001090c00000101ec1b0000040052030000010101fb0e0d0001010101000000010000016c6962726172792f636f72652f7372632f6f7073006c6962726172792f636f72652f7372632f707472006c6962726172792f636f72652f7372632f666d74006c6962726172792f636f72652f737263006c6962726172792f636f72652f7372632f736c6963652f69746572006c6962726172792f636f72652f7372632f697465722f747261697473006c6962726172792f636f72652f7372632f737472006c6962726172792f636f72652f7372632f69746572006c6962726172792f636f72652f7372632f697465722f6164617074657273006c6962726172792f636f72652f7372632f6d656d006c6962726172792f636f72652f7372632f6d6163726f73006c6962726172792f636f72652f7372632f736c696365006c6962726172792f636f72652f7372632f6e756d006c6962726172792f636f72652f7372632f6172726179006c6962726172792f636f72652f7372632f63686172000066756e6374696f6e2e7273000100006d6f642e72730002000072742e72730003000070616e69636b696e672e7273000400006e756d2e727300030000636f6e73745f7074722e727300020000696e7472696e736963732e7273000400006d75745f7074722e7273000200006d6f642e7273000300006d6163726f732e7273000500006974657261746f722e72730006000076616c69646174696f6e732e727300070000616363756d2e727300060000636d702e72730004000072616e67652e7273000800006d61702e72730009000066696c7465722e727300090000636f756e742e727300070000697465722e7273000700006d6f642e7273000a00006f7074696f6e2e7273000400006d6f642e7273000b00006d6f642e727300070000696e6465782e7273000c00007472616974732e7273000700006d6f642e7273000c000075696e745f6d6163726f732e7273000d0000697465722e7273000c0000656e756d65726174652e72730009000063656c6c2e7273000400006275696c646572732e727300030000726573756c742e7273000400006d617962655f756e696e69742e7273000a00006d6f642e7273000e0000636d702e7273000c00007061747465726e2e7273000700006d656d6368722e7273000c00006d6574686f64732e7273000f000000000902a27701000000000003f90101040205090a03860a090000010403050503d375090200010902000001010404000902a677010000000000033301050e0a030f09020001090c000001010402000902b47701000000000003ea030105010a0300090000010902000001010405000902b67701000000000003d2010105170a03130906000106039a7e0918000103e60109040001039a7e0924000105150603e80109020001051e0302090e00010406050d03b505091a00010407050903d20d090200010405051e03fa6c0904000104070509038613090400010406050d03ae72090800010407050903d20d090200010405051503fb6c09080001040705090385130902000106030009040001040505170603f56c0908000106039a7e0906000105140603f901090400010515030209040001051e037f091c000105150302090400010406050d03a305090200010407050903d20d090200010408050d039c73090c00010407050903e40c0902000106038f6b090a000104050514060381020902000105150301090400010408050d038b06090800010405051503f67909020001051e0302090a000105150301090200010406050d039905090400010407050903d20d090200010408050d039c73090c00010407050903e40c0902000106038f6b090800010408050d06038d08090400010405053e03827a09060001050d030209020001050a030109140001060b0300090200010904000001010409000902f87801000000000003dd090105090a03e003091e0001051303a77c090c000106039b76090c000105090603f70d09040001051303ee7b0904000105190305090200010603967609020001050f0603fb090902000105090603000902000103857609040001040a051806038601090200010603fa7e09040001040b05150603b113090400010408050d03dc7409040001040c0505038c7809020001040a051803ed0009080001040d051c03af7f09020001040a051803d100090200010409050d03e50809020001050f031009020001050906030009020001052306030909020001051a06030009040001050906038d0409040001051a03f97b09020001051b03e90009020001053103a47f09060001051503dc000904000106038d7509060001050606039d0a09200001060b0300091c0001050003e3750904000104020509060394090926000106030009060001040905110603f900090400010402050903cd00090a000106030009040001040905110603b37f090400010603f3750914000105090603800b09020001040e05340353090600010409050d032e090400010603ff740910000105150603f30a090200010530030a0904000105230603000904000105300300090200010383750906000105090603800b090c0001040e0534035309040001040f050c039a7a090200010409050d039406090200010603ff74090c000105240603970a090a00010511030109040001030109140001050903fb7e090e0001040e053403bf01090800010409050d03c27e09080001051103fa00091000010603f175091000010603910a090200010301090400010603ee7509080001040e05340603d30a090200010906000001010409000902dc7a01000000000003f2090105140a0301091c0001051103010904000105140302090e0001052c060300090200010b03000912000103897609040001050a0603f80909020001060b0300090a00010904000001010409000902327b01000000000003bb0a01041505120a039b7a090200010409050c03e7050916000104160509039a78090200010409050c03e607090800010518030509040001051d060300090400010406050d0603dc7c09040001040b050903b87b09040001040c05000603a97d09120001041305260603910109040001051106030009020001040b05100603c70109040001040e053403fb0709040001040f050c039a7a09020001040a051803997c09020001040c050d03a07f0904000105080301090800010516030a090400010505035b0904000105110306090400010508032109040001051a0305090400010505035a090400010511060300090200010505030009040001050c06032909040001051e030509040001051203010904000105050351090400010511060300090200010505030009040001050d06032f090400010413050903cb00090200010603f47e09040001040a051806038601091e0001040c050d03a07f090400010508030109040001060359090400010603330908000106034d09040001050c06033b09040001050006034509040001051a060338090400010511035a0904000106030009040001051e06032e09040001051203010904000105050351090400010511060300090600010505030009040001050d06032f090200010413050903cb00090600010417050c03cc000904000105090304090200010418050c037d0904000104170513030f0904000104190509032c090800010603ec7d0904000104150603bc0709020001041903d87a090400010603ec7d0904000104150603bc07090200010603c4780902000104090603d40a0904000105120304090400010412050803c3750908000106036509040001040a051806038601090200010603fa7e09040001040b05150603b113090400010408050d03dc7409040001040c0505038c7809020001040a051803ed0009080001040d051c03af7f09020001040a051803d100090200010402051f03bb0c09040001041a0545036509060001051603800e09080001040a051803e065090600010603fa7e09040001040b05150603b113090200010408050d03dc7409040001040c0505038c7809020001040a051803ed0009080001040d051c03af7f09020001040a051803d100090200010603fa7e090200010386010902000103fa7e09020001040b05150603b113090600010408050d03dc7409040001040c0505038c7809020001040a051803ed0009080001040d051c03af7f09020001040a051803d100090200010603fa7e09020001041205150603c7000922000105000603b97f09060001051b0603fe00090e00010534060300090400010533030009020001051b030009040001041b050d0603e7080902000104120505039a77090400010509035b09020001050c030609020001041c03e80a090200010603b87409020001041a053806039908091200010406050d03867f09040001040a051803e779090600010603fa7e09020001041205190603d0000904000105120301090200010507032309020001050606030009040001051203000902000106035d09020001050503230902000105110360090400010507032009020001050606030009040001051206035d090200010323090200010505060300090200010507030009040001050603000904000105120300090200010505030009020001051206035d0902000105050323090200010511036009020001050703200904000105060603000904000105120300090200010505030009020001040a05180603120904000104120511034e09040001040a05180332090200010603000906000103fa7e090400010386010904000103fa7e09040001038601090600010412051206035d090600010408050d03aa07090200010412050703e7780902000105060603000904000105120300090200010505030009020001040a05180603120904000104120511035e09020001040a05180322090200010603fa7e090400010412051b0603fe00090200010534060300090400010533030009020001051b030009040001041b050d0603e7080902000104120505039a7709040001050d0367090200010409051403f60909020001051b0317090400010535037009060001051503100904000106038d750906000103f30a09260001053006030a0904000105230603000904000105300300090200010383750906000105090603800b090e0001040e0534035309040001040f050c039a7a090200010409050d039406090200010603ff74090c000105280603e30a090a00010515030109040001050903b07e090e0001040e053403bf0109080001040f050c039a7a090400010409050d03a804090400010603eb7609100001040e05340603d30a0902000104090506031609040001060b0300091400010904000001010404000902aa7e01000000000003ed000105050a030709020001090c000001010409000902b87e01000000000003b7080105090a03bb7909180001050b03c90609080001050903b77909040001050503c90609080001050e030e09020001040a051803bc78090400010603fa7e0904000103860109040001040905150603cb0709220001051406030009020001051506030109020001052d0603000904000105150300090400010510060313090600010505060300090200010511060301090200010505060300090400010511060301090400010533036f09020001050503110904000105150304090200010505030f090600010403050c039978090600010603ed7e090a0001051d0603960109040001051b0603000902000103ea7e09020001040905090603eb080902000105190301090400010505030e090800010403050c039978090600010603ed7e090a0001051d0603960109040001051b0603000902000103ea7e09020001040905090603ec0809020001052d0307090400010406050d03ac7e090200010403050903eb7909040001051a060300090200010509030009020001040905110603cc0709040001040a051803b078090200010409051d03b90709100001040a051803c778090400010603fa7e0904000103860109080001040905150603bd0709120001051406030009020001051506030109020001052d060300090400010515030009040001040305090603c67809060001051a060300090200010509030009040001040905110603bc0709040001040a051803c078090200010409051a03d707090a00010418050c03fc78090400010603a77e090600010409051a0603dd08090200010418050c03fc78090400010409051a038407090400010406050d03c27e090400010409050903bf0109040001052106030009040001050903000908000103a2770906000105020603e20809060001060b030009100001090400000101041e000902368001000000000003ba0501040905090a03ba0609000001091200000101041e000902488001000000000003d50501040905090a039f060900000109120000010104200009025a8001000000000003f10c0105050a030109020001090c0000010104150009026880010000000000038a0f01040405050a038b7209020001090c0000010104050009027680010000000000039901010408050d0a03f30609060001040505000603f3770908000106039301090800010421050903d602090200010405051403ea7c090400010603ad7f09080001052306032a0902000103e900090800010603ed7e090400010418050c0603ed03090a00010405050903817d090a0001050e032e09160001060b0300090200010418050d0603d20209040001090e00000101041f000902e680010000000000031e010413050c0a03ce0409460001041a0523039c0d091800010423050d03d26e09040001041f034a090a00010301090400010413050c03c704090e00010424051903b17e090800010418050c0342090a00010425050803cb7d09080001050b030d0906000106034809040001050c0603390902000105090304090c0001050b037b090200010402051f03890d09060001051b03010908000104250508039273090400010603ac7f090e000105100603eb00090600010406050d03b406090400010425051503c679090400010529030409060001041b050d03e508090200010425050503c67609020001051503d2000908000105290304090a0001041b050d03e408090200010425050503c67609020001050903db0009080001050b037209020001050c03580906000105090304090c0001050b037b09020001060348090400010603e1000904000106039f7f09040001050c06033909060001050b037f090c000106034809080001042405200603b403090200010511060300090200010418050c0603ac7f090800010423050d03fb7d090200010424051c03dd02090400010603c87c09040001041f051006032109140001051103010906000106035e090e0001041a050906038912090800010603f76d09040001041f050606032a09100001060b0300091a00010904000001010409000902a28201000000000003a20101052b0a0301090c00010426050803f60b09020001050d031f09040001050f0363090800010513032009060001050d06030009040001051206030109080001050d06030009040001050f060361090c00010513032209060001050d06030009040001051206030109080001050d06030009060001051206030109080001050d060300090400010512060303090c0001050d06030009060001051206030109080001050d06030009060001051206030109080001050d06030009060001051206030109080001050d06030009040001040905090603dc73090a000105060301090a0001060b0300090200010904000001010409000902568301000000000003be010105090a0301090200010506030109300001060b03000902000109040000010104090009028e8301000000000003c5010105090a030109000001090a000001010409000902988301000000000003c9010105090a030109020001052b0359090c00010426050803f60b09020001050d031f09040001050f0363090800010513032009060001050d06030009040001051206030109080001050d06030009040001050f060361090c00010513032209060001050d06030009040001051206030109080001050d06030009060001051206030109080001050d060300090400010512060303090c0001050d06030009060001051206030109080001050d06030009060001051206030109080001050d06030009060001051206030109080001050d06030009040001040905090603dc73090a000105060328090a0001060b03000902000109040000010104090009024e8401000000000003cd010105090a0301090200010371091e00010506031009140001060b030009020001090400000101041f000902888401000000000003b3020105170a0301091200010420050903f10709040001041f03a078090200010603ba7d0908000105100603b602090400010409050903c10b09040001041f050006038972090400010409050903f70d09040001041f05100603bf740904000105000603ca7d09020001051e0603c002090400010603c07d0904000105140603b702090a00010409050903be0909040001041f051503c376091600010603c87d09020001040905090603f50b090e0001041f051e03cb76090a00010409050903b50909020001042003a70309040001041f051103a673090200010409051403e406090c00010603da7609040001041f05210603bb02090200010409051703e806090400010415050903f002090800010409051303947d090a0001051403010904000103010904000105180301090800010509037709080001041f0511039c79091400010409050903e40609040001041f0511039c79090a00010409050903b80909080001041f050006038b740912000105090603b502090200010311090400010506030209060001060b0300091000010904000001010409000902a88501000000000003e40f0105090a03907c090c0001041f050503a376090c00010409050903cf0d090c0001041f050c03fd72090e0001050006039c7d09020001050c03e40209040001039c7d09020001042005090603a60a09020001041f051403c07809020001050006039a7d090a0001051403e60209020001040905090603910b09080001041f051403ef740906000104090509038f0909020001041f051503f2760914000104090509038e0909020001041f03f776091600010409050603fd0c09040001060b0300090a0001090400000101041a0009024086010000000000038a1a01050d0a030109020001090c0000010104090009024e8601000000000003cf110105090a03ec01090000010916000001010422000902648601000000000003820101040905090a03f20a090a00010422051e038f75090200010409050903f10a09020001041f050503a376091000010409050903cf0d090c0001041f050c03fd7209140001050006039c7d09020001050c03e40209040001039c7d09020001042005090603a60a09020001041f051403c07809020001050006039a7d090a0001051403e60209020001040905090603910b09080001041f051403ef740906000104090509038f0909020001041f051503f2760914000104090509038e0909020001041f03f776091600010422050f03977e09040001060b03000908000109040000010104050009020687010000000000039901010408050d0a03f30609060001040505000603f3770908000106039401090800010421050903d502090200010405051403ea7c090400010603ad7f09080001052306032a0902000103ea00090800010603ec7e090400010418050c0603ed03090a00010405050903817d090a0001050e032e09160001060b0300090200010418050d0603d20209040001090e00000101004743433a2028292031322e322e30004c696e6b65723a204c4c442031362e302e32000000000000000000000000000000000000000000000000000000000000010000000400f1ff000000000000000000000000000000000000000000000300fa2601000000000000000000000000000000000000000300fe2601000000000000000000000000000000000000000300322701000000000000000000000000001e00000000000300322701000000000000000000000000002a00000001000500f8bc01000000000010000000000000005300000002000300d6880100000000004c000000000000009b0000000000030030280100000000000000000000000000a70000000100010091040100000000000c00000000000000d30000000000030074280100000000000000000000000000df000000000003009e280100000000000000000000000000eb00000002000300f87401000000000036000000000000004501000002000300c6420100000000000800000000000000540100000200030002950100000000002800000000000000cd010000000003008e290100000000000000000000000000d901000000000300bc290100000000000000000000000000e501000000000300e4290100000000000000000000000000f101000002000300ca7201000000000022000000000000006c020000020003000870010000000000d6000000000000000003000002000300ec720100000000003a000000000000003903000002000300227401000000000042000000000000007803000000000300822a01000000000000000000000000008403000000000300ac2a010000000000000000000000000090030000020003002673010000000000fc000000000000001804000002000300687201000000000062000000000000004b04000000000300f82b0100000000000000000000000000570400000100010056040100000000000c000000000000008204000000000300182c01000000000000000000000000008f040000010001004c040100000000000a00000000000000ba04000002000300fc710100000000006c00000000000000ed040000020003000491010000000000b2000000000000006e05000002000300228d0100000000005400000000000000af05000002000300e88f010000000000a2000000000000004c06000002000300588a0100000000005600000000000000ab06000000000300aa2e0100000000000000000000000000b8060000010001009d040100000000001100000000000000e406000000000300ee2e0100000000000000000000000000f106000000000300182f0100000000000000000000000000fe06000000000300a82f01000000000000000000000000000b07000000000300d62f01000000000000000000000000001807000000000300fe2f010000000000000000000000000025070000000003009c3001000000000000000000000000003207000000000300c63001000000000000000000000000003f0700000200030040860100000000000e00000000000000a50700000000030074320100000000000000000000000000b20700000100010070040100000000002100000000000000bb07000002000300aa7e0100000000000e00000000000000e807000002000300c691010000000000720000000000000069080000020003002a760100000000006001000000000000a508000002000300768d0100000000007c01000000000000eb080000020003008e960100000000007e0500000000000020090000020003002e750100000000007a000000000000006109000002000300fe430100000000005800000000000000b8090000020003004e430100000000005800000000000000140a000002000300a64301000000000058000000000000006e0a00000200030056a30100000000008601000000000000af0a0000020003002a950100000000006401000000000000e90a00000200030052450100000000005800000000000000480b000002000300f6420100000000005800000000000000a30b000002000300249f0100000000009200000000000000de0b000000000300a43b0100000000000000000000000000eb0b00000100010040090100000000001c00000000000000f50b0000000003003e3c0100000000000000000000000000020c00000100010060090100000000002b000000000000002d0c000000000300463c01000000000000000000000000003a0c00000100010018020100000000002000000000000000650c000000000300503c0100000000000000000000000000720c000000000300583c01000000000000000000000000007f0c0000020003005a800100000000000e00000000000000b20c000002000300b69f010000000000a003000000000000f60c000002000300564401000000000052000000000000004f0d000002000300aa450100000000004e00000000000000a20d000002000300a8440100000000005800000000000000f50d00000200030000450100000000005200000000000000550e0000020003000c9c01000000000018030000000000008c0e00000000030024400100000000000000000000000000990e0000000003002c400100000000000000000000000000a60e00000100010090090100000000002000000000000000d10e00000000030072410100000000000000000000000000de0e0000000003007a410100000000000000000000000000eb0e000001000100b0010100000000002000000000000000150f00000000030084410100000000000000000000000000220f0000000003008c4101000000000000000000000000002f0f0000000003009e4101000000000000000000000000003c0f000000000300a6410100000000000000000000000000490f000000000300b0410100000000000000000000000000560f000000000300b8410100000000000000000000000000630f000000000300c2410100000000000000000000000000700f00000100010050070100000000002b000000000000009a0f000000000300d2410100000000000000000000000000a70f000001000100d0010100000000001c00000000000000ad0f000000000300dc410100000000000000000000000000ba0f000001000100f0010100000000002100000000000000c00f000000000300e8410100000000000000000000000000cd0f000000000300f4410100000000000000000000000000da0f00000000030000420100000000000000000000000000000000000000030012420100000000000000000000000000e70f000002000300a6770100000000000e00000000000000181000000200030012420100000000000a000000000000000000000000000300124201000000000000000000000000002a100000020003008a77010000000000180000000000000000000000000003001c4201000000000000000000000000005f100000020003001c420100000000000a0000000000000000000000000003001c4201000000000000000000000000000000000000000300264201000000000000000000000000008a1000000200030026420100000000000a000000000000000000000000000300264201000000000000000000000000000000000000000300304201000000000000000000000000009310000002000300304201000000000008000000000000000000000000000300304201000000000000000000000000009e100000020003004268010000000000d4030000000000000000000000000300384201000000000000000000000000002911000002000300384201000000000008000000000000000000000000000300384201000000000000000000000000003611000002000300166c010000000000f203000000000000000000000000030040420100000000000000000000000000c31100000200030040420100000000004e0000000000000000000000000003004042010000000000000000000000000000000000000003004242010000000000000000000000000000000000000003004c42010000000000000000000000000000000000000003008e420100000000000000000000000000d0110000020003008e42010000000000300000000000000000000000000003008e4201000000000000000000000000000000000000000300904201000000000000000000000000000000000000000300964201000000000000000000000000000000000000000300be420100000000000000000000000000e211000002000300be4201000000000008000000000000000000000000000300be4201000000000000000000000000000000000000000300c64201000000000000000000000000000000000000000300c64201000000000000000000000000000000000000000300ce420100000000000000000000000000ef11000002000300ce4201000000000008000000000000000000000000000300ce4201000000000000000000000000000000000000000300d6420100000000000000000000000000fe11000002000300d64201000000000008000000000000000000000000000300d64201000000000000000000000000000000000000000300de4201000000000000000000000000001212000002000300de420100000000000a000000000000000000000000000300de4201000000000000000000000000000000000000000300e84201000000000000000000000000002d12000002000300e8420100000000000e000000000000000000000000000300e84201000000000000000000000000000000000000000300e84201000000000000000000000000000000000000000300e84201000000000000000000000000000000000000000300ea4201000000000000000000000000000000000000000300ea4201000000000000000000000000000000000000000300ec4201000000000000000000000000000000000000000300f64201000000000000000000000000000000000000000300f64201000000000000000000000000000000000000000300f64201000000000000000000000000000000000000000300f84201000000000000000000000000000000000000000300fc42010000000000000000000000000066120000000003002e43010000000000000000000000000073120000000003003643010000000000000000000000000000000000000003004e43010000000000000000000000000000000000000003004e4301000000000000000000000000000000000000000300504301000000000000000000000000000000000000000300544301000000000000000000000000008012000000000300864301000000000000000000000000008d120000000003008e4301000000000000000000000000000000000000000300a64301000000000000000000000000000000000000000300a64301000000000000000000000000000000000000000300a84301000000000000000000000000000000000000000300ac4301000000000000000000000000009a12000000000300de430100000000000000000000000000a712000000000300e64301000000000000000000000000000000000000000300fe4301000000000000000000000000000000000000000300fe430100000000000000000000000000000000000000030000440100000000000000000000000000000000000000030004440100000000000000000000000000b41200000000030036440100000000000000000000000000c1120000000003003e44010000000000000000000000000000000000000003005644010000000000000000000000000000000000000003005644010000000000000000000000000000000000000003005844010000000000000000000000000000000000000003005a440100000000000000000000000000ce120000020003006a8f0100000000007e000000000000005313000000000300884401000000000000000000000000006013000000000300904401000000000000000000000000000000000000000300a84401000000000000000000000000000000000000000300a84401000000000000000000000000000000000000000300aa4401000000000000000000000000000000000000000300ae4401000000000000000000000000006d13000000000300e04401000000000000000000000000007a13000000000300e84401000000000000000000000000000000000000000300004501000000000000000000000000000000000000000300004501000000000000000000000000000000000000000300024501000000000000000000000000000000000000000300044501000000000000000000000000008713000002000300f28e01000000000078000000000000000d14000000000300324501000000000000000000000000001a140000000003003a45010000000000000000000000000000000000000003005245010000000000000000000000000000000000000003005245010000000000000000000000000000000000000003005445010000000000000000000000000000000000000003005845010000000000000000000000000027140000000003008a4501000000000000000000000000003414000000000300924501000000000000000000000000000000000000000300aa4501000000000000000000000000000000000000000300aa4501000000000000000000000000000000000000000300ac4501000000000000000000000000000000000000000300b04501000000000000000000000000004114000000000300d64501000000000000000000000000004e14000000000300de4501000000000000000000000000000000000000000300f84501000000000000000000000000005b14000002000300f8450100000000009a000000000000000000000000000300f84501000000000000000000000000000000000000000300fa450100000000000000000000000000000000000000030002460100000000000000000000000000a11400000000030018460100000000000000000000000000ae1400000100010038020100000000004000000000000000000000000000030092460100000000000000000000000000ec140000020003009246010000000000dc000000000000000000000000000300924601000000000000000000000000000000000000000300964601000000000000000000000000000000000000000300a24601000000000000000000000000002e150000020003006e47010000000000ee1a00000000000000000000000003006e4701000000000000000000000000007215000000000400e0bb01000000000000000000000000007c15000000000400e8bb01000000000000000000000000008615000000000400f0bb01000000000000000000000000009015000000000400f8bb01000000000000000000000000009a1500000000040000bc0100000000000000000000000000a41500000000040008bc0100000000000000000000000000ae1500000000040010bc0100000000000000000000000000b81500000000040018bc010000000000000000000000000000000000000003006e47010000000000000000000000000000000000000003007047010000000000000000000000000000000000000003008a470100000000000000000000000000c2150000000003000a480100000000000000000000000000cf150000000003001e480100000000000000000000000000dc150000000003006a480100000000000000000000000000e9150000000003007e480100000000000000000000000000f615000000000300c84801000000000000000000000000000316000000000300e24801000000000000000000000000001016000000000300284901000000000000000000000000001d160000000003003e49010000000000000000000000000000000000000003005c6201000000000000000000000000002a160000020003005c62010000000000140400000000000000000000000003005c62010000000000000000000000000000000000000003005e6201000000000000000000000000000000000000000300786201000000000000000000000000006c1600000200030070660100000000003c00000000000000a6160000000003003e630100000000000000000000000000b31600000100010060030100000000001c00000000000000bc16000002000300b6660100000000004c00000000000000f51600000200030002670100000000004c00000000000000401700000200030068800100000000000e000000000000007317000000000300b66501000000000000000000000000008017000000000300ca6501000000000000000000000000008d17000000000300d46501000000000000000000000000009a17000000000300de650100000000000000000000000000a717000000000300e8650100000000000000000000000000b41700000100010000030100000000002100000000000000bd17000000000300f2650100000000000000000000000000ca1700000100010030030100000000002400000000000000d31700000000030000660100000000000000000000000000e0170000000003000a660100000000000000000000000000ed17000001000100d0020100000000002100000000000000f6170000000003001466010000000000000000000000000003180000000003001e6601000000000000000000000000001018000000000300286601000000000000000000000000001d18000001000100a00201000000000023000000000000002618000000000300366601000000000000000000000000003318000001000100a00301000000000010000000000000005e18000000000300506601000000000000000000000000006b18000001000100e80301000000000010000000000000009618000002000300ac660100000000000a00000000000000cc1800000000030062660100000000000000000000000000000000000000030070660100000000000000000000000000000000000000030070660100000000000000000000000000d91800000000030088660100000000000000000000000000e618000000000300966601000000000000000000000000000000000000000300ac6601000000000000000000000000000000000000000300ac6601000000000000000000000000000000000000000300b66601000000000000000000000000000000000000000300b6660100000000000000000000000000f318000000000300d46601000000000000000000000000000019000000000300de6601000000000000000000000000000d19000000000300ec6601000000000000000000000000000000000000000300026701000000000000000000000000000000000000000300026701000000000000000000000000001a190000000003002267010000000000000000000000000027190000000003002c6701000000000000000000000000003419000000000300426701000000000000000000000000004119000001000100f8030100000000000d0000000000000000000000000003004e6701000000000000000000000000006c190000020003004e67010000000000f40000000000000000000000000003004e670100000000000000000000000000ab190000000003001a680100000000000000000000000000b8190000000003002e680100000000000000000000000000c5190000000003003868010000000000000000000000000000000000000003004268010000000000000000000000000000000000000003004268010000000000000000000000000000000000000003004468010000000000000000000000000000000000000003005c680100000000000000000000000000d21900000000030062680100000000000000000000000000df1900000100050050bc010000000000a800000000000000031a0000000003006e680100000000000000000000000000101a000000000300186a01000000000000000000000000001e1a0000000003005a6a01000000000000000000000000002c1a0000000003008a6b01000000000000000000000000003a1a000000000300946b0100000000000000000000000000481a000000000300a26b0100000000000000000000000000561a000000000300b66b0100000000000000000000000000641a000000000300c06b0100000000000000000000000000711a000000000300d46b01000000000000000000000000007e1a000000000300dc6b01000000000000000000000000008c1a00000100010078020100000000002000000000000000b61a000000000300e66b0100000000000000000000000000c31a000000000300ee6b0100000000000000000000000000d01a000000000300f86b0100000000000000000000000000de1a000000000300006c01000000000000000000000000000000000000000300166c01000000000000000000000000000000000000000300166c01000000000000000000000000000000000000000300186c01000000000000000000000000000000000000000300326c0100000000000000000000000000ec1a000000000300326c0100000000000000000000000000fa1a000000000300506c0100000000000000000000000000081b0000000003009c6c0100000000000000000000000000161b000000000300446d0100000000000000000000000000241b000000000300946f0100000000000000000000000000321b0000000003009e6f0100000000000000000000000000401b000000000300ac6f01000000000000000000000000004e1b000000000300c06f01000000000000000000000000005c1b000000000300d86f01000000000000000000000000006a1b000000000300e06f0100000000000000000000000000781b000000000300ea6f0100000000000000000000000000861b000000000300f26f010000000000000000000000000000000000000003000870010000000000000000000000000000000000000003000870010000000000000000000000000000000000000003000a700100000000000000000000000000000000000000030018700100000000000000000000000000941b000002000300de700100000000004a00000000000000dc1b00000200030028710100000000003200000000000000361c000000000300bc700100000000000000000000000000441c000001000100100401000000000019000000000000000000000000000300de7001000000000000000000000000000000000000000300de7001000000000000000000000000000000000000000300e07001000000000000000000000000000000000000000300e470010000000000000000000000000000000000000003002871010000000000000000000000000000000000000003002871010000000000000000000000000000000000000003002a71010000000000000000000000000000000000000003002c7101000000000000000000000000004d1c0000020003005a710100000000006e0000000000000000000000000003005a71010000000000000000000000000000000000000003005a71010000000000000000000000000000000000000003005c710100000000000000000000000000000000000000030062710100000000000000000000000000981c000002000300448801000000000062000000000000000000000000000300c8710100000000000000000000000000cb1c000002000300c87101000000000034000000000000000000000000000300c87101000000000000000000000000000000000000000300ca7101000000000000000000000000000000000000000300cc7101000000000000000000000000000000000000000300fc7101000000000000000000000000000000000000000300fc7101000000000000000000000000000000000000000300fe71010000000000000000000000000000000000000003000a72010000000000000000000000000000000000000003006872010000000000000000000000000000000000000003006872010000000000000000000000000000000000000003006a7201000000000000000000000000000000000000000300767201000000000000000000000000000000000000000300ca7201000000000000000000000000000000000000000300ca7201000000000000000000000000000000000000000300ec7201000000000000000000000000000000000000000300ec7201000000000000000000000000000000000000000300ee7201000000000000000000000000000000000000000300f4720100000000000000000000000000000000000000030026730100000000000000000000000000000000000000030026730100000000000000000000000000000000000000030028730100000000000000000000000000000000000000030036730100000000000000000000000000181d00000000030052730100000000000000000000000000261d00000100010062040100000000000b00000000000000521d000000000300ae730100000000000000000000000000601d000000000300087401000000000000000000000000000000000000000300227401000000000000000000000000000000000000000300227401000000000000000000000000000000000000000300647401000000000000000000000000006e1d00000200030064740100000000009200000000000000000000000000030064740100000000000000000000000000000000000000030066740100000000000000000000000000000000000000030068740100000000000000000000000000c91d0000000003006c740100000000000000000000000000d71d00000000010060010100000000000000000000000000e11d0000000003007a740100000000000000000000000000ea1d00000000030080740100000000000000000000000000f81d0000010001002b050100000000000f00000000000000231e0000000003008c7401000000000000000000000000002c1e000000000300927401000000000000000000000000003a1e00000100010020050100000000000b00000000000000651e0000000003009e7401000000000000000000000000006e1e000000000300a27401000000000000000000000000007c1e000001000100f0040100000000000f00000000000000a71e000000000300aa740100000000000000000000000000b51e00000100010000050100000000002000000000000000e01e000000000300b6740100000000000000000000000000e91e000000000300bc740100000000000000000000000000f71e000000000300cc740100000000000000000000000000001f000000000300d07401000000000000000000000000000e1f000001000100ae040100000000000700000000000000391f000000000300d8740100000000000000000000000000471f000001000100b8040100000000002000000000000000721f000002000300a88501000000000098000000000000000000000000000300f6740100000000000000000000000000b81f000002000300f67401000000000002000000000000000000000000000300f67401000000000000000000000000000000000000000300f87401000000000000000000000000000000000000000300f874010000000000000000000000000000000000000003002e75010000000000000000000000000000000000000003002e7501000000000000000000000000000000000000000300307501000000000000000000000000000000000000000300347501000000000000000000000000000000000000000300a8750100000000000000000000000000f71f000002000300a87501000000000082000000000000000000000000000300a87501000000000000000000000000000000000000000300aa7501000000000000000000000000000000000000000300ae75010000000000000000000000000000000000000003002a76010000000000000000000000000000000000000003002a76010000000000000000000000000000000000000003002e76010000000000000000000000000000000000000003005276010000000000000000000000000000000000000003008a77010000000000000000000000000000000000000003008a7701000000000000000000000000000000000000000300a27701000000000000000000000000003820000002000300a27701000000000004000000000000000000000000000300a27701000000000000000000000000000000000000000300a27701000000000000000000000000000000000000000300a27701000000000000000000000000000000000000000300a27701000000000000000000000000000000000000000300a47701000000000000000000000000000000000000000300a47701000000000000000000000000000000000000000300a67701000000000000000000000000000000000000000300a67701000000000000000000000000000000000000000300a67701000000000000000000000000000000000000000300a67701000000000000000000000000000000000000000300a67701000000000000000000000000000000000000000300a67701000000000000000000000000000000000000000300a87701000000000000000000000000000000000000000300a87701000000000000000000000000000000000000000300aa7701000000000000000000000000000000000000000300b47701000000000000000000000000000000000000000300b47701000000000000000000000000007320000002000300b47701000000000002000000000000000000000000000300b47701000000000000000000000000000000000000000300b47701000000000000000000000000000000000000000300b47701000000000000000000000000000000000000000300b47701000000000000000000000000000000000000000300b67701000000000000000000000000000000000000000300b6770100000000000000000000000000fd2000000000040020bc01000000000000000000000000000721000002000300b67701000000000042010000000000000000000000000300b67701000000000000000000000000000000000000000300b67701000000000000000000000000000000000000000300b67701000000000000000000000000000000000000000300b87701000000000000000000000000000000000000000300ba7701000000000000000000000000000000000000000300bc7701000000000000000000000000003821000000000300c877010000000000000000000000000046210000010001009e05010000000000c8000000000000000000000000000300d47701000000000000000000000000000000000000000300d87701000000000000000000000000007221000000000300dc7701000000000000000000000000000000000000000300fc7701000000000000000000000000000000000000000300fe77010000000000000000000000000000000000000003000c78010000000000000000000000000000000000000003002678010000000000000000000000000000000000000003002678010000000000000000000000000000000000000003002878010000000000000000000000000000000000000003002878010000000000000000000000000000000000000003002c78010000000000000000000000000000000000000003002c78010000000000000000000000000000000000000003003078010000000000000000000000000000000000000003003078010000000000000000000000000000000000000003003878010000000000000000000000000000000000000003003878010000000000000000000000000000000000000003003a78010000000000000000000000000000000000000003003a78010000000000000000000000000000000000000003004278010000000000000000000000000000000000000003004278010000000000000000000000000000000000000003004478010000000000000000000000000000000000000003004478010000000000000000000000000000000000000003004878010000000000000000000000000000000000000003004878010000000000000000000000000000000000000003005078010000000000000000000000000000000000000003005078010000000000000000000000000000000000000003005678010000000000000000000000000000000000000003005a78010000000000000000000000000000000000000003005e78010000000000000000000000000000000000000003007a78010000000000000000000000000000000000000003007e78010000000000000000000000000000000000000003008078010000000000000000000000000000000000000003008078010000000000000000000000000000000000000003008278010000000000000000000000000000000000000003008278010000000000000000000000000000000000000003008e78010000000000000000000000000000000000000003008e78010000000000000000000000000000000000000003009078010000000000000000000000000000000000000003009078010000000000000000000000000000000000000003009a78010000000000000000000000000000000000000003009a78010000000000000000000000000000000000000003009c7801000000000000000000000000000000000000000300a07801000000000000000000000000000000000000000300a87801000000000000000000000000000000000000000300a87801000000000000000000000000000000000000000300aa7801000000000000000000000000000000000000000300aa7801000000000000000000000000000000000000000300b47801000000000000000000000000000000000000000300b67801000000000000000000000000000000000000000300ba7801000000000000000000000000000000000000000300ba7801000000000000000000000000000000000000000300bc7801000000000000000000000000000000000000000300bc7801000000000000000000000000000000000000000300c87801000000000000000000000000000000000000000300c87801000000000000000000000000000000000000000300ca7801000000000000000000000000000000000000000300ca7801000000000000000000000000000000000000000300d27801000000000000000000000000000000000000000300d27801000000000000000000000000000000000000000300d67801000000000000000000000000000000000000000300d67801000000000000000000000000000000000000000300dc7801000000000000000000000000000000000000000300dc7801000000000000000000000000008021000000000300de7801000000000000000000000000008e21000001000100600901000000000000000000000000000000000000000300de780100000000000000000000000000b921000002000300f878010000000000e4010000000000000000000000000300f27801000000000000000000000000000000000000000300f47801000000000000000000000000000000000000000300f87801000000000000000000000000000000000000000300f87801000000000000000000000000000000000000000300f87801000000000000000000000000000000000000000300f87801000000000000000000000000000000000000000300f87801000000000000000000000000000000000000000300fa78010000000000000000000000000000000000000003001479010000000000000000000000000000000000000003001679010000000000000000000000000000000000000003001679010000000000000000000000000000000000000003002279010000000000000000000000000000000000000003002279010000000000000000000000000000000000000003002e79010000000000000000000000000000000000000003003279010000000000000000000000000000000000000003003279010000000000000000000000000000000000000003003679010000000000000000000000000000000000000003003679010000000000000000000000000000000000000003003879010000000000000000000000000000000000000003003a79010000000000000000000000000000000000000003003c79010000000000000000000000000000000000000003003e79010000000000000000000000000000000000000003004279010000000000000000000000000000000000000003004479010000000000000000000000000000000000000003004479010000000000000000000000000000000000000003004879010000000000000000000000000000000000000003004879010000000000000000000000000000000000000003004c79010000000000000000000000000000000000000003005079010000000000000000000000000000000000000003005079010000000000000000000000000000000000000003005279010000000000000000000000000000000000000003005279010000000000000000000000000000000000000003005a79010000000000000000000000000000000000000003005a79010000000000000000000000000000000000000003005c79010000000000000000000000000000000000000003005c79010000000000000000000000000000000000000003005e79010000000000000000000000000000000000000003005e79010000000000000000000000000000000000000003006079010000000000000000000000000000000000000003006079010000000000000000000000000000000000000003006279010000000000000000000000000000000000000003006479010000000000000000000000000000000000000003006679010000000000000000000000000000000000000003006a79010000000000000000000000000000000000000003006e79010000000000000000000000000000000000000003006e79010000000000000000000000000000000000000003007079010000000000000000000000000000000000000003007079010000000000000000000000000000000000000003007279010000000000000000000000000000000000000003007279010000000000000000000000000000000000000003007879010000000000000000000000000000000000000003007879010000000000000000000000000000000000000003007c79010000000000000000000000000000000000000003007c790100000000000000000000000000000000000000030082790100000000000000000000000000000000000000030082790100000000000000000000000000f221000002000300dc7a01000000000056000000000000000000000000000300a27901000000000000000000000000000000000000000300be7901000000000000000000000000000000000000000300c27901000000000000000000000000000000000000000300e87901000000000000000000000000000000000000000300e87901000000000000000000000000000000000000000300ee7901000000000000000000000000000000000000000300ee7901000000000000000000000000000000000000000300f27901000000000000000000000000000000000000000300f27901000000000000000000000000000000000000000300fc7901000000000000000000000000000000000000000300fc7901000000000000000000000000000000000000000300007a01000000000000000000000000000000000000000300007a01000000000000000000000000000000000000000300047a01000000000000000000000000000000000000000300047a01000000000000000000000000000000000000000300187a010000000000000000000000000000000000000003001a7a010000000000000000000000000000000000000003001a7a01000000000000000000000000000000000000000300207a01000000000000000000000000000000000000000300207a01000000000000000000000000000000000000000300247a01000000000000000000000000000000000000000300247a01000000000000000000000000000000000000000300347a01000000000000000000000000000000000000000300347a01000000000000000000000000000000000000000300367a01000000000000000000000000000000000000000300367a010000000000000000000000000000000000000003003a7a010000000000000000000000000000000000000003003e7a01000000000000000000000000000000000000000300407a01000000000000000000000000000000000000000300467a01000000000000000000000000000000000000000300527a01000000000000000000000000000000000000000300567a01000000000000000000000000000000000000000300567a01000000000000000000000000000000000000000300587a01000000000000000000000000000000000000000300587a010000000000000000000000000000000000000003005a7a010000000000000000000000000000000000000003005a7a01000000000000000000000000000000000000000300667a01000000000000000000000000000000000000000300667a01000000000000000000000000000000000000000300707a01000000000000000000000000000000000000000300747a01000000000000000000000000000000000000000300887a01000000000000000000000000000000000000000300967a01000000000000000000000000000000000000000300967a010000000000000000000000000000000000000003009e7a010000000000000000000000000000000000000003009e7a01000000000000000000000000000000000000000300a67a01000000000000000000000000000000000000000300a67a01000000000000000000000000000000000000000300b67a01000000000000000000000000000000000000000300b67a01000000000000000000000000000000000000000300c67a01000000000000000000000000000000000000000300c87a01000000000000000000000000000000000000000300cc7a01000000000000000000000000000000000000000300d47a01000000000000000000000000000000000000000300d67a01000000000000000000000000000000000000000300d67a01000000000000000000000000000000000000000300dc7a01000000000000000000000000000000000000000300dc7a01000000000000000000000000000000000000000300dc7a01000000000000000000000000000000000000000300dc7a01000000000000000000000000000000000000000300dc7a01000000000000000000000000000000000000000300dc7a01000000000000000000000000000000000000000300de7a01000000000000000000000000000000000000000300e87a01000000000000000000000000000000000000000300f87a01000000000000000000000000000000000000000300fc7a010000000000000000000000000000000000000003000a7b010000000000000000000000000000000000000003000c7b010000000000000000000000000000000000000003001e7b01000000000000000000000000000000000000000300227b01000000000000000000000000000000000000000300247b010000000000000000000000000000000000000003002e7b01000000000000000000000000000000000000000300327b01000000000000000000000000000000000000000300327b0100000000000000000000000000392200000000040028bc0100000000000000000000000000432200000000040030bc01000000000000000000000000004d22000002000300327b01000000000078030000000000000000000000000300327b01000000000000000000000000000000000000000300327b01000000000000000000000000000000000000000300327b01000000000000000000000000000000000000000300347b01000000000000000000000000000000000000000300347b01000000000000000000000000000000000000000300347b01000000000000000000000000000000000000000300467b010000000000000000000000000000000000000003004a7b010000000000000000000000000000000000000003004a7b010000000000000000000000000000000000000003004c7b010000000000000000000000000000000000000003004c7b01000000000000000000000000000000000000000300547b01000000000000000000000000000000000000000300547b01000000000000000000000000000000000000000300587b010000000000000000000000000000000000000003005c7b01000000000000000000000000000000000000000300607b01000000000000000000000000000000000000000300607b01000000000000000000000000000000000000000300647b01000000000000000000000000000000000000000300647b01000000000000000000000000000000000000000300767b01000000000000000000000000000000000000000300767b010000000000000000000000000000000000000003007a7b010000000000000000000000000000000000000003007a7b010000000000000000000000000000000000000003007c7b01000000000000000000000000000000000000000300807b01000000000000000000000000000000000000000300807b01000000000000000000000000000000000000000300847b01000000000000000000000000000000000000000300847b01000000000000000000000000000000000000000300867b01000000000000000000000000000000000000000300867b01000000000000000000000000000000000000000300887b01000000000000000000000000000000000000000300887b010000000000000000000000000000000000000003008c7b010000000000000000000000000000000000000003008c7b01000000000000000000000000000000000000000300947b01000000000000000000000000000000000000000300987b010000000000000000000000000000000000000003009c7b010000000000000000000000000000000000000003009c7b01000000000000000000000000000000000000000300a07b01000000000000000000000000000000000000000300a07b01000000000000000000000000000000000000000300a47b01000000000000000000000000000000000000000300a47b01000000000000000000000000000000000000000300a87b01000000000000000000000000000000000000000300ac7b01000000000000000000000000000000000000000300ac7b01000000000000000000000000000000000000000300ae7b01000000000000000000000000000000000000000300b27b01000000000000000000000000000000000000000300b67b01000000000000000000000000000000000000000300b67b01000000000000000000000000000000000000000300ba7b01000000000000000000000000000000000000000300be7b01000000000000000000000000000000000000000300c27b01000000000000000000000000000000000000000300c27b01000000000000000000000000000000000000000300c47b01000000000000000000000000000000000000000300c87b01000000000000000000000000000000000000000300cc7b01000000000000000000000000000000000000000300cc7b01000000000000000000000000000000000000000300ce7b01000000000000000000000000000000000000000300ce7b01000000000000000000000000000000000000000300d27b01000000000000000000000000000000000000000300d27b01000000000000000000000000000000000000000300f07b01000000000000000000000000000000000000000300f07b01000000000000000000000000000000000000000300f47b01000000000000000000000000000000000000000300f47b01000000000000000000000000000000000000000300f87b01000000000000000000000000000000000000000300fc7b01000000000000000000000000000000000000000300047c01000000000000000000000000000000000000000300087c010000000000000000000000000000000000000003000c7c01000000000000000000000000000000000000000300107c01000000000000000000000000000000000000000300147c01000000000000000000000000000000000000000300187c01000000000000000000000000000000000000000300187c010000000000000000000000000000000000000003001c7c010000000000000000000000000000000000000003001c7c01000000000000000000000000000000000000000300207c01000000000000000000000000000000000000000300207c01000000000000000000000000000000000000000300247c01000000000000000000000000000000000000000300287c01000000000000000000000000000000000000000300287c010000000000000000000000000000000000000003002e7c01000000000000000000000000000000000000000300327c01000000000000000000000000000000000000000300347c01000000000000000000000000000000000000000300347c010000000000000000000000000000000000000003003a7c010000000000000000000000000000000000000003003a7c010000000000000000000000000000000000000003003e7c010000000000000000000000000000000000000003003e7c01000000000000000000000000000000000000000300407c01000000000000000000000000000000000000000300447c01000000000000000000000000000000000000000300447c01000000000000000000000000000000000000000300487c01000000000000000000000000000000000000000300487c01000000000000000000000000000000000000000300507c01000000000000000000000000000000000000000300507c01000000000000000000000000000000000000000300547c01000000000000000000000000000000000000000300547c01000000000000000000000000000000000000000300567c01000000000000000000000000000000000000000300567c010000000000000000000000000000000000000003005a7c010000000000000000000000000000000000000003005a7c010000000000000000000000000000000000000003005e7c010000000000000000000000000000000000000003005e7c01000000000000000000000000000000000000000300607c01000000000000000000000000000000000000000300607c01000000000000000000000000000000000000000300627c01000000000000000000000000000000000000000300627c01000000000000000000000000000000000000000300667c010000000000000000000000000000000000000003006a7c01000000000000000000000000000000000000000300727c01000000000000000000000000000000000000000300727c01000000000000000000000000000000000000000300767c01000000000000000000000000000000000000000300787c01000000000000000000000000000000000000000300787c010000000000000000000000000000000000000003007c7c010000000000000000000000000000000000000003007c7c01000000000000000000000000000000000000000300807c01000000000000000000000000000000000000000300847c01000000000000000000000000000000000000000300847c01000000000000000000000000000000000000000300867c01000000000000000000000000000000000000000300867c010000000000000000000000000000000000000003008e7c010000000000000000000000000000000000000003008e7c01000000000000000000000000000000000000000300907c01000000000000000000000000000000000000000300907c01000000000000000000000000000000000000000300927c01000000000000000000000000000000000000000300927c01000000000000000000000000000000000000000300967c01000000000000000000000000000000000000000300967c010000000000000000000000000000000000000003009c7c010000000000000000000000000000000000000003009c7c01000000000000000000000000000000000000000300a47c01000000000000000000000000000000000000000300a47c01000000000000000000000000000000000000000300aa7c01000000000000000000000000000000000000000300aa7c01000000000000000000000000000000000000000300ae7c01000000000000000000000000000000000000000300ae7c01000000000000000000000000000000000000000300b07c01000000000000000000000000000000000000000300b47c01000000000000000000000000000000000000000300b47c01000000000000000000000000000000000000000300b67c01000000000000000000000000000000000000000300b67c01000000000000000000000000000000000000000300be7c01000000000000000000000000000000000000000300be7c01000000000000000000000000000000000000000300c07c01000000000000000000000000000000000000000300c07c01000000000000000000000000000000000000000300c27c01000000000000000000000000000000000000000300c27c01000000000000000000000000000000000000000300c47c01000000000000000000000000000000000000000300c47c01000000000000000000000000000000000000000300c67c01000000000000000000000000000000000000000300c67c01000000000000000000000000000000000000000300c87c01000000000000000000000000000000000000000300c87c01000000000000000000000000000000000000000300ce7c01000000000000000000000000000000000000000300d27c01000000000000000000000000000000000000000300d27c01000000000000000000000000000000000000000300d47c01000000000000000000000000000000000000000300d47c01000000000000000000000000000000000000000300dc7c01000000000000000000000000000000000000000300dc7c01000000000000000000000000000000000000000300de7c01000000000000000000000000000000000000000300de7c01000000000000000000000000000000000000000300e07c01000000000000000000000000000000000000000300e07c01000000000000000000000000000000000000000300e27c01000000000000000000000000000000000000000300e27c01000000000000000000000000007c22000000000300e67c01000000000000000000000000008a22000000000300ee7c01000000000000000000000000000000000000000300047d010000000000000000000000000000000000000003000a7d01000000000000000000000000000000000000000300187d01000000000000000000000000000000000000000300187d010000000000000000000000000000000000000003001c7d010000000000000000000000000000000000000003001e7d01000000000000000000000000000000000000000300227d01000000000000000000000000000000000000000300247d01000000000000000000000000000000000000000300247d01000000000000000000000000000000000000000300287d01000000000000000000000000000000000000000300287d010000000000000000000000000000000000000003002a7d010000000000000000000000000000000000000003002a7d010000000000000000000000000000000000000003002c7d010000000000000000000000000000000000000003002e7d010000000000000000000000000000000000000003002e7d01000000000000000000000000000000000000000300307d010000000000000000000000000000000000000003003a7d010000000000000000000000000000000000000003003e7d01000000000000000000000000000000000000000300427d01000000000000000000000000000000000000000300427d01000000000000000000000000000000000000000300467d01000000000000000000000000000000000000000300467d010000000000000000000000000000000000000003004c7d010000000000000000000000000000000000000003004c7d010000000000000000000000000000000000000003004e7d010000000000000000000000000000000000000003004e7d01000000000000000000000000000000000000000300527d01000000000000000000000000000000000000000300547d01000000000000000000000000000000000000000300567d01000000000000000000000000000000000000000300567d010000000000000000000000000000000000000003005a7d010000000000000000000000000000000000000003005c7d010000000000000000000000000000000000000003005e7d010000000000000000000000000000000000000003005e7d01000000000000000000000000000000000000000300607d01000000000000000000000000000000000000000300607d01000000000000000000000000000000000000000300647d01000000000000000000000000000000000000000300647d01000000000000000000000000000000000000000300667d01000000000000000000000000000000000000000300667d010000000000000000000000000000000000000003006a7d010000000000000000000000000000000000000003006c7d010000000000000000000000000000000000000003006c7d010000000000000000000000000000000000000003006e7d010000000000000000000000000000000000000003006e7d01000000000000000000000000000000000000000300707d01000000000000000000000000000000000000000300747d01000000000000000000000000000000000000000300787d010000000000000000000000000000000000000003007a7d010000000000000000000000000000000000000003007c7d010000000000000000000000000000000000000003007e7d010000000000000000000000000000000000000003007e7d01000000000000000000000000000000000000000300807d01000000000000000000000000000000000000000300807d01000000000000000000000000000000000000000300827d01000000000000000000000000000000000000000300827d01000000000000000000000000000000000000000300867d01000000000000000000000000000000000000000300867d010000000000000000000000000000000000000003008a7d010000000000000000000000000000000000000003008c7d010000000000000000000000000000000000000003008e7d01000000000000000000000000000000000000000300927d01000000000000000000000000000000000000000300927d01000000000000000000000000000000000000000300967d01000000000000000000000000000000000000000300967d01000000000000000000000000000000000000000300987d01000000000000000000000000000000000000000300987d010000000000000000000000000000000000000003009e7d010000000000000000000000000000000000000003009e7d01000000000000000000000000000000000000000300a27d01000000000000000000000000000000000000000300a67d01000000000000000000000000000000000000000300aa7d01000000000000000000000000000000000000000300b07d01000000000000000000000000000000000000000300b67d01000000000000000000000000000000000000000300b67d01000000000000000000000000000000000000000300b87d01000000000000000000000000000000000000000300b87d01000000000000000000000000000000000000000300ba7d01000000000000000000000000000000000000000300ba7d01000000000000000000000000000000000000000300be7d01000000000000000000000000000000000000000300c07d01000000000000000000000000000000000000000300c27d01000000000000000000000000000000000000000300c67d01000000000000000000000000000000000000000300c67d01000000000000000000000000000000000000000300c87d01000000000000000000000000000000000000000300c87d01000000000000000000000000000000000000000300ca7d01000000000000000000000000000000000000000300ca7d01000000000000000000000000000000000000000300ce7d01000000000000000000000000000000000000000300ce7d01000000000000000000000000000000000000000300d07d01000000000000000000000000000000000000000300d07d01000000000000000000000000000000000000000300d47d01000000000000000000000000000000000000000300d67d01000000000000000000000000000000000000000300da7d01000000000000000000000000000000000000000300dc7d01000000000000000000000000000000000000000300dc7d01000000000000000000000000000000000000000300e07d01000000000000000000000000000000000000000300e07d01000000000000000000000000000000000000000300e27d01000000000000000000000000000000000000000300e27d01000000000000000000000000000000000000000300e47d01000000000000000000000000000000000000000300e47d01000000000000000000000000000000000000000300e87d01000000000000000000000000000000000000000300e87d01000000000000000000000000000000000000000300ee7d01000000000000000000000000000000000000000300ee7d01000000000000000000000000000000000000000300f27d01000000000000000000000000000000000000000300f27d01000000000000000000000000000000000000000300f87d01000000000000000000000000000000000000000300f87d010000000000000000000000000000000000000003001e7e010000000000000000000000000000000000000003001e7e01000000000000000000000000000000000000000300227e01000000000000000000000000000000000000000300267e01000000000000000000000000000000000000000300287e010000000000000000000000000000000000000003002e7e010000000000000000000000000000000000000003003c7e01000000000000000000000000000000000000000300407e01000000000000000000000000000000000000000300407e01000000000000000000000000000000000000000300427e01000000000000000000000000000000000000000300427e01000000000000000000000000000000000000000300447e01000000000000000000000000000000000000000300447e01000000000000000000000000000000000000000300507e01000000000000000000000000000000000000000300507e010000000000000000000000000000000000000003005a7e010000000000000000000000000000000000000003005e7e010000000000000000000000000000000000000003006c7e010000000000000000000000000000000000000003006c7e01000000000000000000000000000000000000000300747e01000000000000000000000000000000000000000300747e01000000000000000000000000000000000000000300787e01000000000000000000000000000000000000000300787e010000000000000000000000000000000000000003007c7e010000000000000000000000000000000000000003007c7e010000000000000000000000000000000000000003008c7e010000000000000000000000000000000000000003008e7e010000000000000000000000000000000000000003008e7e01000000000000000000000000000000000000000300927e01000000000000000000000000000000000000000300927e01000000000000000000000000000000000000000300a67e01000000000000000000000000000000000000000300aa7e01000000000000000000000000000000000000000300aa7e01000000000000000000000000000000000000000300aa7e01000000000000000000000000000000000000000300aa7e01000000000000000000000000000000000000000300aa7e01000000000000000000000000000000000000000300ac7e01000000000000000000000000000000000000000300ac7e01000000000000000000000000000000000000000300ae7e01000000000000000000000000000000000000000300b87e01000000000000000000000000000000000000000300b87e01000000000000000000000000009822000002000300b87e0100000000007e010000000000000000000000000300b87e01000000000000000000000000000000000000000300b87e01000000000000000000000000000000000000000300b87e01000000000000000000000000000000000000000300ba7e01000000000000000000000000000000000000000300ca7e01000000000000000000000000000000000000000300d07e01000000000000000000000000000000000000000300d07e01000000000000000000000000000000000000000300d87e01000000000000000000000000000000000000000300d87e01000000000000000000000000000000000000000300dc7e01000000000000000000000000000000000000000300dc7e01000000000000000000000000000000000000000300e47e01000000000000000000000000000000000000000300e47e01000000000000000000000000000000000000000300e67e01000000000000000000000000000000000000000300ea7e01000000000000000000000000000000000000000300ea7e01000000000000000000000000000000000000000300ee7e01000000000000000000000000000000000000000300f27e0100000000000000000000000000bf220000000003000c7f01000000000000000000000000000000000000000300147f01000000000000000000000000000000000000000300147f01000000000000000000000000000000000000000300167f01000000000000000000000000000000000000000300187f010000000000000000000000000000000000000003001c7f01000000000000000000000000000000000000000300207f01000000000000000000000000000000000000000300267f01000000000000000000000000000000000000000300267f01000000000000000000000000000000000000000300287f010000000000000000000000000000000000000003002a7f010000000000000000000000000000000000000003002e7f01000000000000000000000000000000000000000300327f01000000000000000000000000000000000000000300347f01000000000000000000000000000000000000000300347f01000000000000000000000000000000000000000300387f01000000000000000000000000000000000000000300387f010000000000000000000000000000000000000003003a7f01000000000000000000000000000000000000000300407f01000000000000000000000000000000000000000300407f01000000000000000000000000000000000000000300467f01000000000000000000000000000000000000000300467f01000000000000000000000000000000000000000300507f01000000000000000000000000000000000000000300547f01000000000000000000000000000000000000000300567f01000000000000000000000000000000000000000300587f01000000000000000000000000000000000000000300587f010000000000000000000000000000000000000003005a7f010000000000000000000000000000000000000003005e7f01000000000000000000000000000000000000000300667f01000000000000000000000000000000000000000300667f010000000000000000000000000000000000000003006c7f010000000000000000000000000000000000000003006c7f01000000000000000000000000000000000000000300767f010000000000000000000000000000000000000003007a7f010000000000000000000000000000000000000003007c7f010000000000000000000000000000000000000003007e7f010000000000000000000000000000000000000003007e7f01000000000000000000000000000000000000000300807f01000000000000000000000000000000000000000300847f01000000000000000000000000000000000000000300867f01000000000000000000000000000000000000000300867f010000000000000000000000000000000000000003008a7f010000000000000000000000000000000000000003008a7f010000000000000000000000000000000000000003008c7f010000000000000000000000000000000000000003008e7f01000000000000000000000000000000000000000300927f01000000000000000000000000000000000000000300927f01000000000000000000000000000000000000000300947f01000000000000000000000000000000000000000300947f01000000000000000000000000000000000000000300a47f01000000000000000000000000000000000000000300a47f01000000000000000000000000000000000000000300a87f01000000000000000000000000000000000000000300a87f01000000000000000000000000000000000000000300ac7f01000000000000000000000000000000000000000300b47f01000000000000000000000000000000000000000300c67f01000000000000000000000000000000000000000300c67f01000000000000000000000000000000000000000300c87f01000000000000000000000000000000000000000300ca7f01000000000000000000000000000000000000000300ce7f01000000000000000000000000000000000000000300d27f01000000000000000000000000000000000000000300d87f01000000000000000000000000000000000000000300d87f01000000000000000000000000000000000000000300da7f01000000000000000000000000000000000000000300de7f01000000000000000000000000000000000000000300e27f01000000000000000000000000000000000000000300e27f01000000000000000000000000000000000000000300e47f01000000000000000000000000000000000000000300e47f01000000000000000000000000000000000000000300ee7f01000000000000000000000000000000000000000300ee7f01000000000000000000000000000000000000000300f27f01000000000000000000000000000000000000000300f27f01000000000000000000000000000000000000000300f87f01000000000000000000000000000000000000000300f87f01000000000000000000000000000000000000000300fa7f01000000000000000000000000000000000000000300fe7f01000000000000000000000000000000000000000300fe7f010000000000000000000000000000000000000003000280010000000000000000000000000000000000000003000280010000000000000000000000000000000000000003000680010000000000000000000000000000000000000003000680010000000000000000000000000000000000000003000a80010000000000000000000000000000000000000003000a80010000000000000000000000000000000000000003000e80010000000000000000000000000000000000000003001680010000000000000000000000000000000000000003001c800100000000000000000000000000000000000000030022800100000000000000000000000000000000000000030032800100000000000000000000000000000000000000030036800100000000000000000000000000000000000000030036800100000000000000000000000000cd220000020003003680010000000000120000000000000000000000000003003680010000000000000000000000000000000000000003003680010000000000000000000000000000000000000003003680010000000000000000000000000000000000000003003680010000000000000000000000000027230000000003003c80010000000000000000000000000035230000010001003b050100000000000b00000000000000000000000000030048800100000000000000000000000000000000000000030048800100000000000000000000000000000000000000030048800100000000000000000000000000612300000200030048800100000000001200000000000000000000000000030048800100000000000000000000000000000000000000030048800100000000000000000000000000000000000000030048800100000000000000000000000000000000000000030048800100000000000000000000000000be230000000003004e800100000000000000000000000000cc2300000100010046050100000000000e0000000000000000000000000003005a80010000000000000000000000000000000000000003005a80010000000000000000000000000000000000000003005a80010000000000000000000000000000000000000003005a80010000000000000000000000000000000000000003005a80010000000000000000000000000000000000000003005a80010000000000000000000000000000000000000003005c80010000000000000000000000000000000000000003005c80010000000000000000000000000000000000000003005e80010000000000000000000000000000000000000003006880010000000000000000000000000000000000000003006880010000000000000000000000000000000000000003006880010000000000000000000000000000000000000003006880010000000000000000000000000000000000000003006880010000000000000000000000000000000000000003006a80010000000000000000000000000000000000000003006a80010000000000000000000000000000000000000003006a80010000000000000000000000000000000000000003006c800100000000000000000000000000000000000000030076800100000000000000000000000000000000000000030076800100000000000000000000000000000000000000030076800100000000000000000000000000f8230000020003007680010000000000700000000000000000000000000003007680010000000000000000000000000000000000000003007680010000000000000000000000000000000000000003007680010000000000000000000000000000000000000003007880010000000000000000000000000000000000000003007a80010000000000000000000000000000000000000003007c80010000000000000000000000000000000000000003007c80010000000000000000000000000000000000000003008480010000000000000000000000000000000000000003008480010000000000000000000000000000000000000003008c80010000000000000000000000000000000000000003008c80010000000000000000000000000000000000000003008e80010000000000000000000000000000000000000003008e80010000000000000000000000000000000000000003009280010000000000000000000000000000000000000003009280010000000000000000000000000000000000000003009a80010000000000000000000000000000000000000003009c80010000000000000000000000000000000000000003009c8001000000000000000000000000000000000000000300a48001000000000000000000000000000000000000000300a48001000000000000000000000000000000000000000300a88001000000000000000000000000000000000000000300a88001000000000000000000000000000000000000000300b28001000000000000000000000000000000000000000300b28001000000000000000000000000000000000000000300bc8001000000000000000000000000005824000000000300bc80010000000000000000000000000066240000010001009c0501000000000002000000000000000000000000000300bc8001000000000000000000000000000000000000000300d28001000000000000000000000000000000000000000300d28001000000000000000000000000000000000000000300d48001000000000000000000000000000000000000000300d88001000000000000000000000000000000000000000300d88001000000000000000000000000000000000000000300e68001000000000000000000000000000000000000000300e68001000000000000000000000000000000000000000300e6800100000000000000000000000000922400000000040038bc01000000000000000000000000009c2400000000040040bc0100000000000000000000000000a62400000000040048bc0100000000000000000000000000b024000002000300e680010000000000bc010000000000000000000000000300e68001000000000000000000000000000000000000000300e68001000000000000000000000000000000000000000300e68001000000000000000000000000000000000000000300e880010000000000000000000000000000000000000003000281010000000000000000000000000018250000000003000c81010000000000000000000000000026250000000003001481010000000000000000000000000034250000000003001c81010000000000000000000000000000000000000003002c81010000000000000000000000000000000000000003002c81010000000000000000000000000042250000000003003481010000000000000000000000000000000000000003004481010000000000000000000000000000000000000003004481010000000000000000000000000000000000000003004881010000000000000000000000000000000000000003004881010000000000000000000000000000000000000003005281010000000000000000000000000000000000000003005281010000000000000000000000000000000000000003005681010000000000000000000000000000000000000003006481010000000000000000000000000000000000000003006481010000000000000000000000000000000000000003006c81010000000000000000000000000000000000000003006c81010000000000000000000000000000000000000003007681010000000000000000000000000000000000000003007681010000000000000000000000000000000000000003007e81010000000000000000000000000000000000000003007e81010000000000000000000000000000000000000003008481010000000000000000000000000000000000000003008481010000000000000000000000000000000000000003008881010000000000000000000000000000000000000003008a81010000000000000000000000000000000000000003009681010000000000000000000000000000000000000003009881010000000000000000000000000000000000000003009e81010000000000000000000000000000000000000003009e8101000000000000000000000000000000000000000300a68101000000000000000000000000000000000000000300aa8101000000000000000000000000000000000000000300aa8101000000000000000000000000000000000000000300b88101000000000000000000000000000000000000000300be8101000000000000000000000000000000000000000300c28101000000000000000000000000000000000000000300c28101000000000000000000000000000000000000000300c68101000000000000000000000000000000000000000300c68101000000000000000000000000000000000000000300cc8101000000000000000000000000000000000000000300ce8101000000000000000000000000000000000000000300ce8101000000000000000000000000000000000000000300d08101000000000000000000000000000000000000000300d08101000000000000000000000000000000000000000300d88101000000000000000000000000000000000000000300d88101000000000000000000000000000000000000000300e28101000000000000000000000000000000000000000300e48101000000000000000000000000000000000000000300e48101000000000000000000000000000000000000000300e68101000000000000000000000000000000000000000300e68101000000000000000000000000000000000000000300ee8101000000000000000000000000000000000000000300ee8101000000000000000000000000000000000000000300f08101000000000000000000000000000000000000000300f68101000000000000000000000000000000000000000300f681010000000000000000000000000000000000000003000282010000000000000000000000000000000000000003000482010000000000000000000000000000000000000003000882010000000000000000000000000000000000000003000882010000000000000000000000000000000000000003000c82010000000000000000000000000000000000000003001082010000000000000000000000000000000000000003001682010000000000000000000000000000000000000003001682010000000000000000000000000000000000000003002282010000000000000000000000000000000000000003002a82010000000000000000000000000000000000000003002a82010000000000000000000000000000000000000003002c82010000000000000000000000000000000000000003002e82010000000000000000000000000000000000000003003682010000000000000000000000000000000000000003003682010000000000000000000000000000000000000003003882010000000000000000000000000000000000000003003882010000000000000000000000000000000000000003003c82010000000000000000000000000000000000000003003c82010000000000000000000000000000000000000003004082010000000000000000000000000000000000000003004082010000000000000000000000000000000000000003005482010000000000000000000000000000000000000003005a82010000000000000000000000000000000000000003006882010000000000000000000000000000000000000003007082010000000000000000000000000000000000000003007082010000000000000000000000000000000000000003007482010000000000000000000000000000000000000003007482010000000000000000000000000000000000000003008482010000000000000000000000000000000000000003009e8201000000000000000000000000000000000000000300a28201000000000000000000000000000000000000000300a28201000000000000000000000000005025000002000300a282010000000000b4000000000000000000000000000300a28201000000000000000000000000000000000000000300a28201000000000000000000000000000000000000000300a28201000000000000000000000000000000000000000300a48201000000000000000000000000000000000000000300a68201000000000000000000000000000000000000000300ae8201000000000000000000000000000000000000000300b08201000000000000000000000000000000000000000300b08201000000000000000000000000000000000000000300b48201000000000000000000000000000000000000000300b48201000000000000000000000000000000000000000300bc8201000000000000000000000000000000000000000300bc8201000000000000000000000000000000000000000300c28201000000000000000000000000000000000000000300c28201000000000000000000000000000000000000000300c68201000000000000000000000000000000000000000300ce8201000000000000000000000000000000000000000300d28201000000000000000000000000000000000000000300de8201000000000000000000000000000000000000000300de8201000000000000000000000000000000000000000300e48201000000000000000000000000000000000000000300e48201000000000000000000000000000000000000000300e88201000000000000000000000000000000000000000300f08201000000000000000000000000000000000000000300f68201000000000000000000000000000000000000000300fe82010000000000000000000000000000000000000003000283010000000000000000000000000000000000000003000e83010000000000000000000000000000000000000003001483010000000000000000000000000000000000000003001c83010000000000000000000000000000000000000003002283010000000000000000000000000000000000000003002a83010000000000000000000000000000000000000003003083010000000000000000000000000000000000000003003883010000000000000000000000000000000000000003003c83010000000000000000000000000000000000000003004683010000000000000000000000000000000000000003004683010000000000000000000000000000000000000003005083010000000000000000000000000000000000000003005283010000000000000000000000000000000000000003005683010000000000000000000000000000000000000003005683010000000000000000000000000083250000020003005683010000000000380000000000000000000000000003005683010000000000000000000000000000000000000003005683010000000000000000000000000000000000000003005683010000000000000000000000000000000000000003005883010000000000000000000000000000000000000003005883010000000000000000000000000000000000000003005a830100000000000000000000000000b42500000000030074830100000000000000000000000000c2250000010001006806010000000000300000000000000000000000000003008883010000000000000000000000000000000000000003008a83010000000000000000000000000000000000000003008e83010000000000000000000000000000000000000003008e830100000000000000000000000000ee250000020003008e830100000000000a0000000000000000000000000003008e83010000000000000000000000000000000000000003008e83010000000000000000000000000000000000000003008e83010000000000000000000000000000000000000003008e83010000000000000000000000000000000000000003009883010000000000000000000000000000000000000003009883010000000000000000000000000044260000020003009883010000000000b60000000000000000000000000003009883010000000000000000000000000000000000000003009883010000000000000000000000000000000000000003009883010000000000000000000000000000000000000003009a83010000000000000000000000000000000000000003009a83010000000000000000000000000000000000000003009c8301000000000000000000000000000000000000000300a68301000000000000000000000000000000000000000300a68301000000000000000000000000000000000000000300a88301000000000000000000000000000000000000000300a88301000000000000000000000000000000000000000300ac8301000000000000000000000000000000000000000300ac8301000000000000000000000000000000000000000300b48301000000000000000000000000000000000000000300b48301000000000000000000000000000000000000000300ba8301000000000000000000000000000000000000000300ba8301000000000000000000000000000000000000000300be8301000000000000000000000000000000000000000300c68301000000000000000000000000000000000000000300ca8301000000000000000000000000000000000000000300d68301000000000000000000000000000000000000000300d68301000000000000000000000000000000000000000300dc8301000000000000000000000000000000000000000300dc8301000000000000000000000000000000000000000300e08301000000000000000000000000000000000000000300e88301000000000000000000000000000000000000000300ee8301000000000000000000000000000000000000000300f68301000000000000000000000000000000000000000300fa83010000000000000000000000000000000000000003000684010000000000000000000000000000000000000003000c84010000000000000000000000000000000000000003001484010000000000000000000000000000000000000003001a84010000000000000000000000000000000000000003002284010000000000000000000000000000000000000003002884010000000000000000000000000000000000000003003084010000000000000000000000000000000000000003003484010000000000000000000000000000000000000003003e84010000000000000000000000000000000000000003003e84010000000000000000000000000000000000000003004884010000000000000000000000000000000000000003004884010000000000000000000000000000000000000003004a84010000000000000000000000000000000000000003004e84010000000000000000000000000000000000000003004e8401000000000000000000000000009c260000020003004e840100000000003a0000000000000000000000000003004e84010000000000000000000000000000000000000003004e84010000000000000000000000000000000000000003004e840100000000000000000000000000000000000000030050840100000000000000000000000000000000000000030050840100000000000000000000000000000000000000030052840100000000000000000000000000f2260000000003006e84010000000000000000000000000000000000000003006e84010000000000000000000000000000000000000003006e84010000000000000000000000000000000000000003008284010000000000000000000000000000000000000003008284010000000000000000000000000000000000000003008484010000000000000000000000000000000000000003008884010000000000000000000000000000000000000003008884010000000000000000000000000000270000020003008884010000000000200100000000000000000000000003008884010000000000000000000000000000000000000003008884010000000000000000000000000000000000000003008884010000000000000000000000000000000000000003008a84010000000000000000000000000000000000000003009884010000000000000000000000000000000000000003009a84010000000000000000000000000000000000000003009e84010000000000000000000000000000000000000003009e8401000000000000000000000000000000000000000300a08401000000000000000000000000000000000000000300a08401000000000000000000000000000000000000000300a88401000000000000000000000000000000000000000300ac8401000000000000000000000000000000000000000300ac8401000000000000000000000000000000000000000300b08401000000000000000000000000000000000000000300b08401000000000000000000000000000000000000000300b48401000000000000000000000000000000000000000300b48401000000000000000000000000000000000000000300b88401000000000000000000000000000000000000000300b88401000000000000000000000000000000000000000300bc8401000000000000000000000000000000000000000300bc8401000000000000000000000000000000000000000300be8401000000000000000000000000000000000000000300c28401000000000000000000000000003c27000000000300c68401000000000000000000000000004a27000001000100960501000000000002000000000000000000000000000300c68401000000000000000000000000000000000000000300d08401000000000000000000000000000000000000000300d48401000000000000000000000000000000000000000300d48401000000000000000000000000007627000000000300de8401000000000000000000000000008427000001000100980501000000000002000000000000000000000000000300ea8401000000000000000000000000000000000000000300ea8401000000000000000000000000000000000000000300ec840100000000000000000000000000b027000000000300f2840100000000000000000000000000be270000010001009a0501000000000001000000000000000000000000000300fa8401000000000000000000000000000000000000000300fa84010000000000000000000000000000000000000003000485010000000000000000000000000000000000000003000485010000000000000000000000000000000000000003000685010000000000000000000000000000000000000003000685010000000000000000000000000000000000000003000a85010000000000000000000000000000000000000003000a85010000000000000000000000000000000000000003000c85010000000000000000000000000000000000000003000c85010000000000000000000000000000000000000003001885010000000000000000000000000000000000000003001885010000000000000000000000000000000000000003001c85010000000000000000000000000000000000000003001c85010000000000000000000000000000000000000003001e85010000000000000000000000000000000000000003002285010000000000000000000000000000000000000003002285010000000000000000000000000000000000000003002a85010000000000000000000000000000000000000003002a85010000000000000000000000000000000000000003003485010000000000000000000000000000000000000003003485010000000000000000000000000000000000000003003885010000000000000000000000000000000000000003003c85010000000000000000000000000000000000000003004485010000000000000000000000000000000000000003004c850100000000000000000000000000000000000000030060850100000000000000000000000000000000000000030060850100000000000000000000000000000000000000030064850100000000000000000000000000ea2700000000030064850100000000000000000000000000f8270000010001005805010000000000300000000000000000000000000003006485010000000000000000000000000000000000000003006e85010000000000000000000000000000000000000003006e85010000000000000000000000000000000000000003007685010000000000000000000000000000000000000003007685010000000000000000000000000024280000000003007c85010000000000000000000000000032280000010001009405010000000000020000000000000000000000000003008885010000000000000000000000000000000000000003008885010000000000000000000000000000000000000003008a85010000000000000000000000000000000000000003008a85010000000000000000000000000000000000000003008e8501000000000000000000000000000000000000000300948501000000000000000000000000000000000000000300a48501000000000000000000000000000000000000000300a88501000000000000000000000000000000000000000300a88501000000000000000000000000000000000000000300a88501000000000000000000000000000000000000000300a88501000000000000000000000000000000000000000300a88501000000000000000000000000000000000000000300aa8501000000000000000000000000000000000000000300b28501000000000000000000000000000000000000000300b48501000000000000000000000000000000000000000300b48501000000000000000000000000000000000000000300c08501000000000000000000000000000000000000000300c08501000000000000000000000000000000000000000300cc8501000000000000000000000000000000000000000300cc8501000000000000000000000000000000000000000300da8501000000000000000000000000000000000000000300da8501000000000000000000000000000000000000000300dc8501000000000000000000000000000000000000000300e08501000000000000000000000000000000000000000300e28501000000000000000000000000000000000000000300e48501000000000000000000000000000000000000000300e48501000000000000000000000000000000000000000300e68501000000000000000000000000000000000000000300e68501000000000000000000000000000000000000000300f08501000000000000000000000000000000000000000300f28501000000000000000000000000000000000000000300fa8501000000000000000000000000000000000000000300fa8501000000000000000000000000000000000000000300008601000000000000000000000000000000000000000300008601000000000000000000000000000000000000000300028601000000000000000000000000000000000000000300028601000000000000000000000000005e28000000000300088601000000000000000000000000006c280000010001009b05010000000000010000000000000000000000000003001686010000000000000000000000000000000000000003001686010000000000000000000000000000000000000003001886010000000000000000000000000000000000000003001886010000000000000000000000000098280000000003001e860100000000000000000000000000a6280000010001003a05010000000000010000000000000000000000000003002e86010000000000000000000000000000000000000003002e86010000000000000000000000000000000000000003003286010000000000000000000000000000000000000003003286010000000000000000000000000000000000000003003c86010000000000000000000000000000000000000003004086010000000000000000000000000000000000000003004086010000000000000000000000000000000000000003004086010000000000000000000000000000000000000003004086010000000000000000000000000000000000000003004086010000000000000000000000000000000000000003004286010000000000000000000000000000000000000003004286010000000000000000000000000000000000000003004486010000000000000000000000000000000000000003004e86010000000000000000000000000000000000000003004e860100000000000000000000000000d2280000020003004e86010000000000160000000000000000000000000003004e86010000000000000000000000000000000000000003004e8601000000000000000000000000001a290000000003004e86010000000000000000000000000000000000000003004e86010000000000000000000000000028290000010001009806010000000000020000000000000000000000000003004e86010000000000000000000000000000000000000003006486010000000000000000000000000000000000000003006486010000000000000000000000000000000000000003006486010000000000000000000000000054290000020003006486010000000000a20000000000000000000000000003006486010000000000000000000000000000000000000003006486010000000000000000000000000000000000000003006486010000000000000000000000000000000000000003006686010000000000000000000000000000000000000003006c86010000000000000000000000000000000000000003006e86010000000000000000000000000000000000000003006e860100000000000000000000000000000000000000030070860100000000000000000000000000000000000000030070860100000000000000000000000000000000000000030072860100000000000000000000000000000000000000030072860100000000000000000000000000b52900000000030076860100000000000000000000000000c329000001000100c006010000000000110000000000000000000000000003008286010000000000000000000000000000000000000003008286010000000000000000000000000000000000000003008e860100000000000000000000000000ef290000000003008e860100000000000000000000000000fd29000001000100a006010000000000200000000000000000000000000003008e8601000000000000000000000000000000000000000300a28601000000000000000000000000000000000000000300a28601000000000000000000000000000000000000000300a48601000000000000000000000000000000000000000300a88601000000000000000000000000000000000000000300aa8601000000000000000000000000000000000000000300ac8601000000000000000000000000000000000000000300ac8601000000000000000000000000000000000000000300ae8601000000000000000000000000000000000000000300ae8601000000000000000000000000000000000000000300b88601000000000000000000000000000000000000000300ba8601000000000000000000000000000000000000000300c28601000000000000000000000000000000000000000300c28601000000000000000000000000000000000000000300c88601000000000000000000000000000000000000000300c88601000000000000000000000000000000000000000300ca8601000000000000000000000000000000000000000300ca860100000000000000000000000000292a000000000300d08601000000000000000000000000000000000000000300de8601000000000000000000000000000000000000000300de8601000000000000000000000000000000000000000300e08601000000000000000000000000000000000000000300e0860100000000000000000000000000372a000000000300e68601000000000000000000000000000000000000000300f68601000000000000000000000000000000000000000300f68601000000000000000000000000000000000000000300fa8601000000000000000000000000000000000000000300fa860100000000000000000000000000000000000000030002870100000000000000000000000000000000000000030006870100000000000000000000000000000000000000030006870100000000000000000000000000452a0000020003000687010000000000700000000000000000000000000003000687010000000000000000000000000000000000000003000687010000000000000000000000000000000000000003000687010000000000000000000000000000000000000003000887010000000000000000000000000000000000000003000a87010000000000000000000000000000000000000003000c87010000000000000000000000000000000000000003000c87010000000000000000000000000000000000000003001487010000000000000000000000000000000000000003001487010000000000000000000000000000000000000003001c87010000000000000000000000000000000000000003001c87010000000000000000000000000000000000000003001e87010000000000000000000000000000000000000003001e87010000000000000000000000000000000000000003002287010000000000000000000000000000000000000003002287010000000000000000000000000000000000000003002a87010000000000000000000000000000000000000003002c87010000000000000000000000000000000000000003002c87010000000000000000000000000000000000000003003487010000000000000000000000000000000000000003003487010000000000000000000000000000000000000003003887010000000000000000000000000000000000000003003887010000000000000000000000000000000000000003004287010000000000000000000000000000000000000003004287010000000000000000000000000000000000000003004c870100000000000000000000000000a52a0000000003004c87010000000000000000000000000000000000000003004c870100000000000000000000000000000000000000030062870100000000000000000000000000000000000000030062870100000000000000000000000000000000000000030064870100000000000000000000000000000000000000030068870100000000000000000000000000000000000000030068870100000000000000000000000000000000000000030076870100000000000000000000000000000000000000030076870100000000000000000000000000000000000000030076870100000000000000000000000000b32a000002000300768701000000000052000000000000000000000000000300768701000000000000000000000000000000000000000300788701000000000000000000000000000000000000000300828701000000000000000000000000005f2b000002000300c8870100000000007c000000000000000000000000000300c88701000000000000000000000000000000000000000300c88701000000000000000000000000000000000000000300ca8701000000000000000000000000000000000000000300d087010000000000000000000000000000000000000003004488010000000000000000000000000000000000000003004488010000000000000000000000000000000000000003004688010000000000000000000000000000000000000003004e8801000000000000000000000000000000000000000300a6880100000000000000000000000000b92b000002000300a68801000000000030000000000000000000000000000300a68801000000000000000000000000000000000000000300d68801000000000000000000000000000000000000000300d68801000000000000000000000000000000000000000300d88801000000000000000000000000000000000000000300dc880100000000000000000000000000000000000000030022890100000000000000000000000000012c0000020003002289010000000000680000000000000000000000000003002289010000000000000000000000000000000000000003002489010000000000000000000000000000000000000003002e890100000000000000000000000000422c0000020003008a890100000000007c0000000000000000000000000003008a89010000000000000000000000000000000000000003008a89010000000000000000000000000000000000000003008c8901000000000000000000000000000000000000000300928901000000000000000000000000009c2c000002000300068a01000000000052000000000000000000000000000300068a01000000000000000000000000000000000000000300068a01000000000000000000000000000000000000000300088a010000000000000000000000000000000000000003000e8a01000000000000000000000000000000000000000300588a01000000000000000000000000000000000000000300588a010000000000000000000000000000000000000003005a8a010000000000000000000000000000000000000003005e8a01000000000000000000000000000000000000000300ae8a0100000000000000000000000000cf2c000002000300ae8a01000000000082010000000000000000000000000300ae8a01000000000000000000000000000000000000000300b08a01000000000000000000000000000000000000000300be8a0100000000000000000000000000002d000000000300908b01000000000000000000000000000e2d000001000100a0070100000000001c00000000000000182d0000000003009a8b0100000000000000000000000000262d000000000300a48b0100000000000000000000000000342d000000000300b88b0100000000000000000000000000422d000000000300c08b0100000000000000000000000000502d000001000100f80601000000000020000000000000007a2d000000000300ce8b0100000000000000000000000000882d00000100010006080100000000002f00000000000000b32d000000000300dc8b0100000000000000000000000000c12d00000100010035080100000000003200000000000000ec2d000000000300f68b0100000000000000000000000000fa2d000000000300fe8b0100000000000000000000000000082e00000100010080070100000000002000000000000000322e000000000300188c0100000000000000000000000000402e000001000100bc070100000000001c000000000000006b2e000000000300228c0100000000000000000000000000792e000001000100d8070100000000002e000000000000000000000000000300308c0100000000000000000000000000a42e000002000300308c01000000000028000000000000000000000000000300308c0100000000000000000000000000ff2e000000000300368c01000000000000000000000000000d2f000001000100280a0100000000005000000000000000772f000000000300408c0100000000000000000000000000852f000001000100780a01000000000050000000000000000000000000000300588c0100000000000000000000000000f32f000002000300588c01000000000062000000000000000000000000000300588c010000000000000000000000000000000000000003005a8c01000000000000000000000000002c300000000003007a8c01000000000000000000000000003a30000000000300868c010000000000000000000000000048300000010001001807010000000000180000000000000072300000000003008e8c0100000000000000000000000000803000000100010030070100000000002000000000000000aa30000000000300a48c0100000000000000000000000000b830000001000100670801000000000026000000000000000000000000000300ba8c0100000000000000000000000000e330000002000300ba8c01000000000068000000000000000000000000000300ba8c01000000000000000000000000000000000000000300bc8c01000000000000000000000000000000000000000300c08c01000000000000000000000000002231000000000300ec8c01000000000000000000000000003031000000000300f48c01000000000000000000000000003e310000000003000e8d01000000000000000000000000004c310000010001008d080100000000000d000000000000000000000000000300228d01000000000000000000000000000000000000000300228d01000000000000000000000000000000000000000300248d01000000000000000000000000000000000000000300288d01000000000000000000000000007731000000000300608d01000000000000000000000000000000000000000300768d01000000000000000000000000000000000000000300768d01000000000000000000000000000000000000000300788d010000000000000000000000000000000000000003008a8d01000000000000000000000000008531000000000300108e010000000000000000000000000093310000000003009e8e0100000000000000000000000000a131000000000300a88e0100000000000000000000000000af310000010001009a080100000000000e00000000000000da31000000000300b48e0100000000000000000000000000e831000000000300be8e0100000000000000000000000000f631000000000300c88e01000000000000000000000000000432000000000300d28e01000000000000000000000000001232000000000300dc8e01000000000000000000000000000000000000000300f28e01000000000000000000000000000000000000000300f28e01000000000000000000000000000000000000000300f48e01000000000000000000000000000000000000000300fa8e01000000000000000000000000002032000000000300348f01000000000000000000000000002e320000000003003c8f01000000000000000000000000003c32000000000300568f01000000000000000000000000004a32000001000100a8080100000000000e0000000000000000000000000003006a8f010000000000000000000000000000000000000003006a8f010000000000000000000000000000000000000003006c8f01000000000000000000000000000000000000000300728f01000000000000000000000000007532000000000300b28f01000000000000000000000000008332000000000300ba8f01000000000000000000000000009132000000000300d48f01000000000000000000000000009f32000001000100b6080100000000000d000000000000000000000000000300e88f01000000000000000000000000000000000000000300e88f01000000000000000000000000000000000000000300ea8f01000000000000000000000000000000000000000300f28f0100000000000000000000000000ca3200000000030054900100000000000000000000000000d8320000000003005c900100000000000000000000000000e63200000000030076900100000000000000000000000000f432000001000100c308010000000000120000000000000000000000000003008a9001000000000000000000000000001f330000020003008a900100000000007a0000000000000000000000000003008a90010000000000000000000000000000000000000003008c9001000000000000000000000000000000000000000300929001000000000000000000000000008333000000000300e290010000000000000000000000000000000000000003000491010000000000000000000000000000000000000003000491010000000000000000000000000000000000000003000691010000000000000000000000000000000000000003001291010000000000000000000000000091330000000003006c9101000000000000000000000000009f33000001000100d80801000000000020000000000000000000000000000300b6910100000000000000000000000000ca33000002000300b69101000000000010000000000000000000000000000300b69101000000000000000000000000000000000000000300c69101000000000000000000000000000000000000000300c69101000000000000000000000000000000000000000300c89101000000000000000000000000000000000000000300d09101000000000000000000000000001b340000000003001a92010000000000000000000000000000000000000003003892010000000000000000000000000029340000020003003892010000000000ca0200000000000000000000000003003892010000000000000000000000000000000000000003003a92010000000000000000000000000000000000000003004a920100000000000000000000000000b334000000000300c4940100000000000000000000000000c134000000000300d8940100000000000000000000000000cf34000000000300e2940100000000000000000000000000dd34000000000300ea940100000000000000000000000000000000000000030002950100000000000000000000000000000000000000030002950100000000000000000000000000eb3400000000030004950100000000000000000000000000f934000000000100880101000000000000000000000000000435000000000300149501000000000000000000000000000e350000000003001695010000000000000000000000000018350000000003001895010000000000000000000000000022350000000003001c9501000000000000000000000000002c350000000003002095010000000000000000000000000000000000000003002a95010000000000000000000000000000000000000003002a95010000000000000000000000000000000000000003002c95010000000000000000000000000000000000000003003c95010000000000000000000000000000000000000003008e96010000000000000000000000000000000000000003008e9601000000000000000000000000000000000000000300929601000000000000000000000000000000000000000300b69601000000000000000000000000003635000000000300169a01000000000000000000000000004435000000000300989b0100000000000000000000000000523500000100010030040100000000001c000000000000005b35000000000300a29b01000000000000000000000000006935000000000300ac9b01000000000000000000000000007735000000000300b69b01000000000000000000000000008535000000000300c09b01000000000000000000000000009335000000000300de9b0100000000000000000000000000a135000000000300e69b0100000000000000000000000000af35000001000100b009010000000000200000000000000000000000000003000c9c010000000000000000000000000000000000000003000c9c010000000000000000000000000000000000000003000e9c01000000000000000000000000000000000000000300249c0100000000000000000000000000da35000000000300e29e0100000000000000000000000000e835000000000300f69e0100000000000000000000000000f635000001000100d0090100000000002b000000000000002236000000000300049f010000000000000000000000000030360000000003000c9f01000000000000000000000000000000000000000300249f01000000000000000000000000000000000000000300249f01000000000000000000000000000000000000000300269f010000000000000000000000000000000000000003002c9f01000000000000000000000000000000000000000300b69f01000000000000000000000000000000000000000300b69f01000000000000000000000000000000000000000300b89f01000000000000000000000000000000000000000300d29f01000000000000000000000000003e360000000003000aa301000000000000000000000000004c360000000003001ea301000000000000000000000000005a3600000000030026a3010000000000000000000000000068360000000003003ea301000000000000000000000000007636000001000100fb090100000000002900000000000000000000000000030056a30100000000000000000000000000000000000000030056a30100000000000000000000000000000000000000030058a30100000000000000000000000000000000000000030064a30100000000000000000000000000a236000000000300b6a401000000000000000000000000000000000000000300dca40100000000000000000000000000b03600000100060008bd0100000000000010080000000000db3600000100060008cd09000000000000100000000000000c370000010001007c0301000000000023000000000000003737000001000100b00301000000000033000000000000006237000001000100f8080100000000000a000000000000008d3700000100010002090100000000000a00000000000000b8370000010001000c090100000000000b00000000000000e337000001000100170901000000000006000000000000000e380000010001001d09010000000000060000000000000039380000010001002309010000000000090000000000000064380000010001002c0901000000000006000000000000000000000000000800000000000000000000000000000000000000000000000b00962900000000000000000000000000000000000000000b00d44200000000000000000000000000008f38000000000f00000000000000000000000000000000000000000000000b002c1200000000000000000000000000000000000000000b00452d00000000000000000000000000000000000000000b00000000000000000000000000000000000000000000000b00914b00000000000000000000000000000000000000000b00643500000000000000000000000000000000000000000800510000000000000000000000000000000000000000000b0020160000000000000000000000000000a338000000000f005c0000000000000000000000000000000000000000000a00700e00000000000000000000000000000000000000000b00011900000000000000000000000000000000000000000b001f0500000000000000000000000000000000000000000b007d0c00000000000000000000000000000000000000000b00561600000000000000000000000000000000000000000b00dc3200000000000000000000000000000000000000000b002b0c00000000000000000000000000000000000000000b00323c00000000000000000000000000000000000000000b00973000000000000000000000000000000000000000000b00e63500000000000000000000000000000000000000000b00982300000000000000000000000000000000000000000b00c52800000000000000000000000000000000000000000b00ec2100000000000000000000000000000000000000000b000c2b00000000000000000000000000000000000000000b00dc4500000000000000000000000000000000000000000b00573800000000000000000000000000000000000000000b006f3700000000000000000000000000000000000000000b00c50b00000000000000000000000000000000000000000b00f90300000000000000000000000000000000000000000b00ad0c00000000000000000000000000000000000000000b00353f00000000000000000000000000000000000000000b00b03000000000000000000000000000000000000000000b00531700000000000000000000000000000000000000000b004d0b00000000000000000000000000000000000000000b00d53400000000000000000000000000000000000000000b00a60000000000000000000000000000000000000000000b00844600000000000000000000000000000000000000000b00fe1200000000000000000000000000000000000000000b00de4000000000000000000000000000000000000000000b002f4500000000000000000000000000000000000000000b002b0500000000000000000000000000000000000000000b00060800000000000000000000000000000000000000000b00cc0000000000000000000000000000000000000000000b00362800000000000000000000000000000000000000000b00933000000000000000000000000000000000000000000b005c1200000000000000000000000000000000000000000b00903100000000000000000000000000000000000000000b00124800000000000000000000000000000000000000000b00752700000000000000000000000000000000000000000b00023e00000000000000000000000000000000000000000b00371300000000000000000000000000000000000000000b00d34500000000000000000000000000000000000000000b002c3b00000000000000000000000000000000000000000b00694800000000000000000000000000000000000000000b008a2e00000000000000000000000000000000000000000b00c21500000000000000000000000000000000000000000b00763500000000000000000000000000000000000000000a00000000000000000000000000000000000000000000000a00400000000000000000000000000000000000000000000a00700000000000000000000000000000000000000000000a00a00000000000000000000000000000000000000000000b00a30b00000000000000000000000000000000000000000b00682b00000000000000000000000000000000000000000b005d3b00000000000000000000000000000000000000000b00e52d00000000000000000000000000000000000000000b006f2900000000000000000000000000000000000000000b004b2900000000000000000000000000000000000000000b00021400000000000000000000000000000000000000000b00d81b00000000000000000000000000000000000000000b00ff4300000000000000000000000000000000000000000b00d04600000000000000000000000000000000000000000b00ba3800000000000000000000000000000000000000000b00771400000000000000000000000000000000000000000b002a2e00000000000000000000000000000000000000000a00200900000000000000000000000000000000000000000a00500900000000000000000000000000000000000000000a00800900000000000000000000000000000000000000000a00b00900000000000000000000000000000000000000000a00e00900000000000000000000000000000000000000000b00650700000000000000000000000000000000000000000b00733200000000000000000000000000000000000000000b006f0700000000000000000000000000000000000000000b001f0300000000000000000000000000000000000000000a00800d00000000000000000000000000000000000000000a00b00d00000000000000000000000000000000000000000a00e00d00000000000000000000000000000000000000000a00100e00000000000000000000000000000000000000000a00400e00000000000000000000000000000000000000000b00ec4900000000000000000000000000000000000000000b00370a00000000000000000000000000000000000000000b006c0a00000000000000000000000000000000000000000b007f0300000000000000000000000000000000000000000b008e2e00000000000000000000000000000000000000000b00de4800000000000000000000000000000000000000000b00ca4000000000000000000000000000000000000000000b00b90c00000000000000000000000000000000000000000b00230500000000000000000000000000000000000000000b00890200000000000000000000000000000000000000000b00cc3100000000000000000000000000000000000000000a00d00000000000000000000000000000000000000000000a00100100000000000000000000000000000000000000000a00400100000000000000000000000000000000000000000a00700100000000000000000000000000000000000000000a00a00100000000000000000000000000000000000000000a00d00100000000000000000000000000000000000000000a00000200000000000000000000000000000000000000000a00300200000000000000000000000000000000000000000a00800200000000000000000000000000000000000000000b008d4700000000000000000000000000000000000000000b00202e00000000000000000000000000000000000000000a00b00200000000000000000000000000000000000000000a00e00200000000000000000000000000000000000000000a00100300000000000000000000000000000000000000000a00400300000000000000000000000000000000000000000a00700300000000000000000000000000000000000000000a00a00300000000000000000000000000000000000000000a00d00300000000000000000000000000000000000000000a00000400000000000000000000000000000000000000000a00300400000000000000000000000000000000000000000a00800400000000000000000000000000000000000000000a00b00400000000000000000000000000000000000000000a00000500000000000000000000000000000000000000000a00300500000000000000000000000000000000000000000a00800500000000000000000000000000000000000000000a00b00500000000000000000000000000000000000000000a00f00500000000000000000000000000000000000000000a00600600000000000000000000000000000000000000000a00b00600000000000000000000000000000000000000000a00f00600000000000000000000000000000000000000000a00200700000000000000000000000000000000000000000a00500700000000000000000000000000000000000000000b00283800000000000000000000000000000000000000000b00d52d00000000000000000000000000000000000000000b005e1700000000000000000000000000000000000000000b005e2b00000000000000000000000000000000000000000b00123100000000000000000000000000000000000000000b003e2900000000000000000000000000000000000000000b00412700000000000000000000000000000000000000000b006a1c00000000000000000000000000000000000000000b001f0700000000000000000000000000000000000000000b007e2300000000000000000000000000000000000000000b00451a00000000000000000000000000000000000000000b001f1700000000000000000000000000000000000000000b00222f00000000000000000000000000000000000000000b00282f00000000000000000000000000000000000000000b009c4900000000000000000000000000000000000000000b00ff1900000000000000000000000000000000000000000b00fa0800000000000000000000000000000000000000000b00584900000000000000000000000000000000000000000b00420f00000000000000000000000000000000000000000b001f0900000000000000000000000000000000000000000b00313900000000000000000000000000000000000000000a00800700000000000000000000000000000000000000000a00b00700000000000000000000000000000000000000000a00e00700000000000000000000000000000000000000000a00100800000000000000000000000000000000000000000a00400800000000000000000000000000000000000000000a00700800000000000000000000000000000000000000000a00a00800000000000000000000000000000000000000000a00e00800000000000000000000000000000000000000000b00f10100000000000000000000000000000000000000000b00ab3c00000000000000000000000000000000000000000b00a93800000000000000000000000000000000000000000b00d83700000000000000000000000000000000000000000b007e3500000000000000000000000000000000000000000a00100a00000000000000000000000000000000000000000a00400a00000000000000000000000000000000000000000a00700a00000000000000000000000000000000000000000a00a00a00000000000000000000000000000000000000000a00d00a00000000000000000000000000000000000000000a00000b00000000000000000000000000000000000000000b00383d00000000000000000000000000000000000000000b00b94400000000000000000000000000000000000000000b00920400000000000000000000000000000000000000000b00f81900000000000000000000000000000000000000000b00232300000000000000000000000000000000000000000b00642900000000000000000000000000000000000000000b005c4900000000000000000000000000000000000000000b00714600000000000000000000000000000000000000000b00bd0900000000000000000000000000000000000000000a00b00b00000000000000000000000000000000000000000a00e00b00000000000000000000000000000000000000000a00100c00000000000000000000000000000000000000000a00400c00000000000000000000000000000000000000000a00700c00000000000000000000000000000000000000000a00b00c00000000000000000000000000000000000000000b00e41c00000000000000000000000000000000000000000b00784700000000000000000000000000000000000000000b00a91c00000000000000000000000000000000000000000b00e02d00000000000000000000000000000000000000000b00f10800000000000000000000000000000000000000000b000b3500000000000000000000000000000000000000000b00553100000000000000000000000000000000000000000b00132300000000000000000000000000000000000000000b000f3000000000000000000000000000000000000000000a00300b00000000000000000000000000000000000000000b00741800000000000000000000000000000000000000000b00153000000000000000000000000000000000000000000b00884400000000000000000000000000000000000000000b00664b00000000000000000000000000000000000000000b00bc4700000000000000000000000000000000000000000b00eb4100000000000000000000000000000000000000000b00164200000000000000000000000000000000000000000a00700b00000000000000000000000000000000000000000b00823700000000000000000000000000000000000000000b00780900000000000000000000000000000000000000000b00db0f00000000000000000000000000000000000000000b00210c00000000000000000000000000000000000000000b004b3000000000000000000000000000000000000000000b00261000000000000000000000000000000000000000000b00783900000000000000000000000000000000000000000b00e34900000000000000000000000000000000000000000b00624800000000000000000000000000000000000000000b00820900000000000000000000000000000000000000000b00ca4b00000000000000000000000000000000000000000b00812700000000000000000000000000000000000000000b001d0e00000000000000000000000000000000000000000b00834700000000000000000000000000000000000000000b00f31500000000000000000000000000000000000000000b00242e00000000000000000000000000000000000000000b00e73c00000000000000000000000000000000000000000b000a1200000000000000000000000000000000000000000b006c0f00000000000000000000000000000000000000000b004b3100000000000000000000000000000000000000000b007c3900000000000000000000000000000000000000000b00f90900000000000000000000000000000000000000000b008f1000000000000000000000000000000000000000000b009d3100000000000000000000000000000000000000000b00211d00000000000000000000000000000000000000000b00a02300000000000000000000000000000000000000000b00663300000000000000000000000000000000000000000b00194500000000000000000000000000000000000000000b00b23a00000000000000000000000000000000000000000b00c10100000000000000000000000000000000000000000b00922a00000000000000000000000000000000000000000b00fd4000000000000000000000000000000000000000000b00804a00000000000000000000000000000000000000000b00e13d00000000000000000000000000000000000000000b00201b00000000000000000000000000000000000000000b008d3c00000000000000000000000000000000000000000b00383600000000000000000000000000000000000000000b00120000000000000000000000000000000000000000000b00241a00000000000000000000000000000000000000000b00522d00000000000000000000000000000000000000000b001e4900000000000000000000000000000000000000000b00e13100000000000000000000000000000000000000000b00fc2100000000000000000000000000000000000000000b000c2200000000000000000000000000000000000000000b004b3400000000000000000000000000000000000000000b00764a00000000000000000000000000000000000000000b00ef3600000000000000000000000000000000000000000b00c20a00000000000000000000000000000000000000000b009c3a00000000000000000000000000000000000000000b009b0b00000000000000000000000000000000000000000b009a1b00000000000000000000000000000000000000000b00b34100000000000000000000000000000000000000000b008b1100000000000000000000000000000000000000000b00511a00000000000000000000000000000000000000000b00d01a00000000000000000000000000000000000000000b00272800000000000000000000000000000000000000000b00b44300000000000000000000000000000000000000000b00a54600000000000000000000000000000000000000000b00ac2500000000000000000000000000000000000000000b00823d00000000000000000000000000000000000000000b00b30500000000000000000000000000000000000000000b00993d00000000000000000000000000000000000000000b00194100000000000000000000000000000000000000000b00b00800000000000000000000000000000000000000000b00652800000000000000000000000000000000000000000b00b12800000000000000000000000000000000000000000b00e13700000000000000000000000000000000000000000b008b3a00000000000000000000000000000000000000000b007a1900000000000000000000000000000000000000000b00d21100000000000000000000000000000000000000000b006d4100000000000000000000000000000000000000000b006a2f00000000000000000000000000000000000000000b00462600000000000000000000000000000000000000000b00280900000000000000000000000000000000000000000b00a90d00000000000000000000000000000000000000000b00f11700000000000000000000000000000000000000000b004c0400000000000000000000000000000000000000000b00d01900000000000000000000000000000000000000000b000f0700000000000000000000000000000000000000000b006e4200000000000000000000000000000000000000000b00663900000000000000000000000000000000000000000b00b40300000000000000000000000000000000000000000b004a0500000000000000000000000000000000000000000b00d93100000000000000000000000000000000000000000b00613400000000000000000000000000000000000000000b00172900000000000000000000000000000000000000000b00400d00000000000000000000000000000000000000000b00001200000000000000000000000000000000000000000b000b3e00000000000000000000000000000000000000000b00fe3000000000000000000000000000000000000000000b00793700000000000000000000000000000000000000000b00fa0100000000000000000000000000000000000000000b00f94500000000000000000000000000000000000000000b007b2f00000000000000000000000000000000000000000b00931700000000000000000000000000000000000000000b00ea1400000000000000000000000000000000000000000b00ec0c00000000000000000000000000000000000000000b00264900000000000000000000000000000000000000000b00811400000000000000000000000000000000000000000b00843b00000000000000000000000000000000000000000b00de1b00000000000000000000000000000000000000000b002d3d00000000000000000000000000000000000000000b00d92d00000000000000000000000000000000000000000b00ff1700000000000000000000000000000000000000000b00923b00000000000000000000000000000000000000000b00ca3b00000000000000000000000000000000000000000b00374700000000000000000000000000000000000000000b005b1c00000000000000000000000000000000000000000b009d0f00000000000000000000000000000000000000000b007f3e00000000000000000000000000000000000000000b004b2d00000000000000000000000000000000000000000b00d72900000000000000000000000000000000000000000b000c4300000000000000000000000000000000000000000b005f1200000000000000000000000000000000000000000b00ab2300000000000000000000000000000000000000000b003c3c00000000000000000000000000000000000000000b00833f00000000000000000000000000000000000000000b007b3600000000000000000000000000000000000000000b00f60000000000000000000000000000000000000000000b003a0800000000000000000000000000000000000000000b00e10e00000000000000000000000000000000000000000b00a71000000000000000000000000000000000000000000b00ad1000000000000000000000000000000000000000000b008b2700000000000000000000000000000000000000000b00873900000000000000000000000000000000000000000b00b50c00000000000000000000000000000000000000000b00564000000000000000000000000000000000000000000b00b71000000000000000000000000000000000000000000b007b4600000000000000000000000000000000000000000b00982e00000000000000000000000000000000000000000b009c2e00000000000000000000000000000000000000000b00261d00000000000000000000000000000000000000000b00fd4900000000000000000000000000000000000000000b00214300000000000000000000000000000000000000000b00431f00000000000000000000000000000000000000000b00f64900000000000000000000000000000000000000000b00790700000000000000000000000000000000000000000b009f1200000000000000000000000000000000000000000b000c0000000000000000000000000000000000000000000b00224500000000000000000000000000000000000000000b006b1600000000000000000000000000000000000000000b00590000000000000000000000000000000000000000000b00161b00000000000000000000000000000000000000000b00fe0500000000000000000000000000000000000000000b00022600000000000000000000000000000000000000000b006d1300000000000000000000000000000000000000000b00532200000000000000000000000000000000000000000b002d0800000000000000000000000000000000000000000b00564500000000000000000000000000000000000000000b00f12000000000000000000000000000000000000000000b008f4600000000000000000000000000000000000000000b00022100000000000000000000000000000000000000000b00080000000000000000000000000000000000000000000b00760a00000000000000000000000000000000000000000b000c1a00000000000000000000000000000000000000000b004e0e00000000000000000000000000000000000000000b00154300000000000000000000000000000000000000000b00e51e00000000000000000000000000000000000000000b00790800000000000000000000000000000000000000000b006b1900000000000000000000000000000000000000000b00a63d00000000000000000000000000000000000000000b00241300000000000000000000000000000000000000000b004b2a00000000000000000000000000000000000000000b00d20100000000000000000000000000000000000000000b006d4800000000000000000000000000000000000000000b00064a00000000000000000000000000000000000000000b001f0100000000000000000000000000000000000000000b005a1a00000000000000000000000000000000000000000b00f62f00000000000000000000000000000000000000000b00972600000000000000000000000000000000000000000b00b00b00000000000000000000000000000000000000000b00e14100000000000000000000000000000000000000000b00092c00000000000000000000000000000000000000000b00043000000000000000000000000000000000000000000b00b60a00000000000000000000000000000000000000000b00413d00000000000000000000000000000000000000000b007b3c00000000000000000000000000000000000000000b00e02900000000000000000000000000000000000000000b00c23600000000000000000000000000000000000000000b00030f00000000000000000000000000000000000000000b001f2a00000000000000000000000000000000000000000b00972100000000000000000000000000000000000000000b00d92100000000000000000000000000000000000000000b003d3600000000000000000000000000000000000000000b00e33300000000000000000000000000000000000000000b00e12700000000000000000000000000000000000000000b00984600000000000000000000000000000000000000000b00f60c00000000000000000000000000000000000000000b002f2a00000000000000000000000000000000000000000b00e93300000000000000000000000000000000000000000b00253400000000000000000000000000000000000000000b000a0400000000000000000000000000000000000000000b001d3d00000000000000000000000000000000000000000b00a73000000000000000000000000000000000000000000b00240100000000000000000000000000000000000000000b00460500000000000000000000000000000000000000000b00224700000000000000000000000000000000000000000b00fa4a00000000000000000000000000000000000000000b002a4700000000000000000000000000000000000000000b00e52600000000000000000000000000000000000000000b008b2c00000000000000000000000000000000000000000b00263200000000000000000000000000000000000000000b002b4500000000000000000000000000000000000000000b00533a00000000000000000000000000000000000000000b00371a00000000000000000000000000000000000000000b00a33100000000000000000000000000000000000000000b00820e00000000000000000000000000000000000000000b00a32b00000000000000000000000000000000000000000b006b1400000000000000000000000000000000000000000b00314400000000000000000000000000000000000000000b00c64600000000000000000000000000000000000000000b00f00c00000000000000000000000000000000000000000b00ec0000000000000000000000000000000000000000000b00061900000000000000000000000000000000000000000b00e03300000000000000000000000000000000000000000b000a2300000000000000000000000000000000000000000b00c03800000000000000000000000000000000000000000b00552900000000000000000000000000000000000000000b00094400000000000000000000000000000000000000000b00312f00000000000000000000000000000000000000000b006b3700000000000000000000000000000000000000000b002f4900000000000000000000000000000000000000000b00402a00000000000000000000000000000000000000000b00cc0800000000000000000000000000000000000000000b00330800000000000000000000000000000000000000000b00a03000000000000000000000000000000000000000000b00a40e00000000000000000000000000000000000000000b00370500000000000000000000000000000000000000000b00774300000000000000000000000000000000000000000b007c3a00000000000000000000000000000000000000000b00ba0300000000000000000000000000000000000000000b00094100000000000000000000000000000000000000000b00910600000000000000000000000000000000000000000b00f50d00000000000000000000000000000000000000000b00023f00000000000000000000000000000000000000000b00583900000000000000000000000000000000000000000b008d2d00000000000000000000000000000000000000000b00b94600000000000000000000000000000000000000000b00294600000000000000000000000000000000000000000b00594b00000000000000000000000000000000000000000b00cb1900000000000000000000000000000000000000000b003c2600000000000000000000000000000000000000000b00bf4400000000000000000000000000000000000000000b001c3200000000000000000000000000000000000000000b00c20200000000000000000000000000000000000000000b00fb1300000000000000000000000000000000000000000b00ec0400000000000000000000000000000000000000000b001e1200000000000000000000000000000000000000000b00714700000000000000000000000000000000000000000b00313200000000000000000000000000000000000000000b00a71800000000000000000000000000000000000000000b00cd0600000000000000000000000000000000000000000b00d73b00000000000000000000000000000000000000000b00413000000000000000000000000000000000000000000b00923e00000000000000000000000000000000000000000b005b0900000000000000000000000000000000000000000b00912600000000000000000000000000000000000000000b00e71700000000000000000000000000000000000000000b008a2200000000000000000000000000000000000000000b00b02b00000000000000000000000000000000000000000b002e1000000000000000000000000000000000000000000a00f00c00000000000000000000000000000000000000000a00200d00000000000000000000000000000000000000000a00500d00000000000000000000000000000000000000000b008c0600000000000000000000000000000000000000000b00033500000000000000000000000000000000000000000b00022d00000000000000000000000000000000000000000b00301800000000000000000000000000000000000000000b00391800000000000000000000000000000000000000000b00352d00000000000000000000000000000000000000000b00731500000000000000000000000000000000000000000b007c4400000000000000000000000000000000000000000300f64201000000000000000000000000000000000000000300a67701000000000000000000000000000000000000000300b47701000000000000000000000000000000000000000300b67701000000000000000000000000000000000000000300f87801000000000000000000000000000000000000000300dc7a01000000000000000000000000000000000000000300327b01000000000000000000000000000000000000000300aa7e01000000000000000000000000000000000000000300b87e010000000000000000000000000000000000000003003680010000000000000000000000000000000000000003004880010000000000000000000000000000000000000003005a8001000000000000000000000000000000000000000300688001000000000000000000000000000000000000000300768001000000000000000000000000000000000000000300e68001000000000000000000000000000000000000000300a282010000000000000000000000000000000000000003005683010000000000000000000000000000000000000003008e83010000000000000000000000000000000000000003009883010000000000000000000000000000000000000003004e8401000000000000000000000000000000000000000300888401000000000000000000000000000000000000000300a885010000000000000000000000000000000000000003004086010000000000000000000000000000000000000003004e860100000000000000000000000000000000000000030064860100000000000000000000000000000000000000030006870100000000000000000000000000000000000000030076870100000000000000000000000000b73800000400f1ff00000000000000000000000000000000bd38000000000300dca40100000000000000000000000000c038000000000300aaa50100000000000000000000000000c338000000000300d2a90100000000000000000000000000c638000000000300f8a90100000000000000000000000000c938000000000300a8a50100000000000000000000000000cd3800000000030098a50100000000000000000000000000d138000000000300cea90100000000000000000000000000d63800000000030086a60100000000000000000000000000db38000000000300cea50100000000000000000000000000e03800000000030070a80100000000000000000000000000e538000000000300caa50100000000000000000000000000ea380000000003009aa60100000000000000000000000000ef3800000000030046a60100000000000000000000000000f43800000000030004a60100000000000000000000000000f93800000000030008a90100000000000000000000000000fe3800000000030014a6010000000000000000000000000003390000000003006ca60100000000000000000000000000083900000000030078a601000000000000000000000000000d390000000003005aa8010000000000000000000000000012390000000003004ea70100000000000000000000000000173900000000030038a901000000000000000000000000001c390000000003007aa801000000000000000000000000002139000000000300e4a601000000000000000000000000002639000000000300e8a701000000000000000000000000002b3900000000030030a80100000000000000000000000000303900000000030056a8010000000000000000000000000035390000000003007ca601000000000000000000000000003a390000000003009ca801000000000000000000000000003f3900000000030012a90100000000000000000000000000443900000000030062a901000000000000000000000000004939000000000300e2a501000000000000000000000000004e39000000000300e8a901000000000000000000000000005439000000000300eca901000000000000000000000000005a39000000000300d4a901000000000000000000000000006039000000000300d8aa01000000000000000000000000006639000000000300b8ab01000000000000000000000000006c39000000000300dcaa0100000000000000000000000000723900000000030044ab01000000000000000000000000007839000000000300beab01000000000000000000000000007e39000000000300baab010000000000000000000000000084390000000003005aaa01000000000000000000000000008a390000000003002eab01000000000000000000000000009039000000000300d4ab01000000000000000000000000009639000000000300faaa01000000000000000000000000009c39000000000300f4aa0100000000000000000000000000a239000000000300c4ab0100000000000000000000000000a83900000000030018ab0100000000000000000000000000ae39000000000300d8ab0100000000000000000000000000b4390000000003005cab0100000000000000000000000000ba3900000000030056ab0100000000000000000000000000c039000000000300c8ab0100000000000000000000000000c63900000000030084ab0100000000000000000000000000cc39000000000300a6ab0100000000000000000000000000d239000000000300a4ab0100000000000000000000000000d839000000000300a0ab0100000000000000000000000000de390000000003000eab0100000000000000000000000000e4390000000003006eab0100000000000000000000000000003a000002020300dca4010000000000ce00000000000000073a000002020300aaa501000000000028040000000000000e3a000002020300d2a90100000000002600000000000000153a000002020300f8a9010000000000e601000000000000ea39000012000300fa26010000000000181b000000000000f939000010000300e4260100000000000000000000000000002e726f64617461002e65685f6672616d65002e74657874002e7364617461002e64617461002e627373002e64656275675f616262726576002e64656275675f696e666f002e64656275675f6172616e676573002e64656275675f72616e676573002e64656275675f737472002e64656275675f7075626e616d6573002e64656275675f7075627479706573002e72697363762e61747472696275746573002e64656275675f6c696e65002e636f6d6d656e74002e73796d746162002e7368737472746162002e73747274616200007374616b652e333936663965326636373736336630382d6367752e30002e4c706372656c5f686930005f5a4e37636b625f73746433656e7634415247563137683861626337373932303633656163623745005f5a4e35616c6c6f63377261775f7665633139526177566563244c54245424432441244754243131616c6c6f636174655f696e3137683961373435623837316432623838663945002e4c706372656c5f686931002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e343330002e4c706372656c5f686933002e4c706372656c5f686932005f5a4e34636f726533707472353564726f705f696e5f706c616365244c54246d6f6c6563756c652e2e6572726f722e2e566572696669636174696f6e4572726f72244754243137683733613437386435323862633430643345005f5f727573745f6465616c6c6f63005f5a4e39305f244c54247574696c2e2e6572726f722e2e4572726f72247532302461732475323024636f72652e2e636f6e766572742e2e46726f6d244c5424636b625f7374642e2e6572726f722e2e5379734572726f7224475424244754243466726f6d3137683035613866363565623361306264316345002e4c706372656c5f686934002e4c706372656c5f686935002e4c706372656c5f686936005f5a4e34636f726535736c69636535696e64657837345f244c5424696d706c2475323024636f72652e2e6f70732e2e696e6465782e2e496e646578244c542449244754242475323024666f72247532302424753562245424753564242447542435696e6465783137683064326565363561653136626361336545005f5a4e3131315f244c5424616c6c6f632e2e7665632e2e566563244c54245424475424247532302461732475323024616c6c6f632e2e7665632e2e737065635f66726f6d5f697465725f6e65737465642e2e5370656346726f6d497465724e6573746564244c5424542443244924475424244754243966726f6d5f697465723137683032353562336632346332623633633445005f5a4e35616c6c6f63337665633136566563244c542454244324412447542434707573683137683832346530366138613965323339383745005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f7233616e793137683031323866356465313834336464653445002e4c706372656c5f686938002e4c706372656c5f686937005f5a4e3130325f244c5424636b625f7374616e64616c6f6e655f74797065732e2e67656e6572617465642e2e626c6f636b636861696e2e2e42797465735265616465722475323024617324753230246d6f6c6563756c652e2e7072656c7564652e2e52656164657224475424367665726966793137683135663233383466353032373265326345005f5a4e386d6f6c6563756c6535627974657335427974657335736c6963653137683339643866386561613338343133646245002e4c706372656c5f686939002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e3936002e4c706372656c5f68693130002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e3234005f5a4e386d6f6c6563756c6535627974657335427974657335736c6963653137683133633337653065643765643238336345005f5a4e39385f244c54246d6f6c6563756c65322e2e7265616465722e2e437572736f72247532302461732475323024636f72652e2e636f6e766572742e2e46726f6d244c5424616c6c6f632e2e7665632e2e566563244c542475382447542424475424244754243466726f6d3137686365383937663564613837343036643045005f5a4e396d6f6c6563756c65323672656164657236437572736f723135736c6963655f62795f6f66667365743137683635646335653064333235363034343945005f5a4e396d6f6c6563756c6532367265616465723130385f244c5424696d706c2475323024636f72652e2e636f6e766572742e2e46726f6d244c54246d6f6c6563756c65322e2e7265616465722e2e437572736f72244754242475323024666f722475323024616c6c6f632e2e7665632e2e566563244c5424753824475424244754243466726f6d3137683965653331373661666261663535343545005f5a4e36345f244c5424616c6c6f632e2e72632e2e5263244c54245424475424247532302461732475323024636f72652e2e6f70732e2e64726f702e2e44726f70244754243464726f703137683663346239333364656266363135663545002e4c706372656c5f68693136002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e383436002e4c706372656c5f68693138002e4c706372656c5f68693137002e4c706372656c5f68693139002e4c706372656c5f68693230002e4c706372656c5f68693231002e4c706372656c5f68693233002e4c706372656c5f68693232005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243135636f70795f66726f6d5f736c69636531376c656e5f6d69736d617463685f6661696c3137686531663934356265353831313135613845002e4c706372656c5f68693131007374722e342e3436005f5a4e34636f72653970616e69636b696e673570616e69633137686437373538656430613265383739363145005f5a4e39385f244c5424636b625f7374642e2e686967685f6c6576656c2e2e517565727949746572244c54244624475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683764366161393561356131323831396645005f5a4e37636b625f7374643130686967685f6c6576656c31346c6f61645f63656c6c5f646174613137683061353964663134343334336539316145005f5a4e396d6f6c6563756c65323672656164657236437572736f7232307461626c655f736c6963655f62795f696e6465783137686232343839353738643638326165663045005f5a4e347574696c3668656c70657231356765745f7363726970745f686173683137686133663334636563626161396538326445005f5a4e37636b625f7374643130686967685f6c6576656c31396c6f61645f63656c6c5f6c6f636b5f686173683137683339633636646239366138646337393445005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f72656164657237547970654964733134787564745f747970655f686173683137686334653636633566343738343237356145005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f726561646572375479706549647331397374616b655f736d745f636f64655f686173683137683939313230643232643561376161363745005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f726561646572375479706549647331377374616b655f736d745f747970655f69643137683133613730383736373561386135323245005f5a4e347574696c3668656c70657232376765745f63656c6c5f636f756e745f62795f747970655f686173683137683433316433366633633236643131663045005f5a4e347574696c3668656c7065723230636865636b5f787564745f747970655f686173683137683030353064373537353834646533643045005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231355374616b65417443656c6c4461746131366d657461646174615f747970655f69643137683136353731366261626264366365656645005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f72656164657237547970654964733138636865636b706f696e745f747970655f69643137683062376537323033303666383865346345005f5a4e347574696c3668656c70657232316765745f787564745f62795f747970655f686173683137686230346631613436386437663535383945002e4c706372656c5f68693238007374722e302e333134002e4c706372656c5f68693132002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e3436002e4c706372656c5f68693133002e4c616e6f6e2e30656130363565396135373639326336653434396165616266643062303633332e3139002e4c706372656c5f68693134002e4c706372656c5f68693135005f5a4e34636f726536726573756c743133756e777261705f6661696c65643137683030653934303161326339653536633045005f5a4e347574696c3668656c70657233306765745f7374616b655f61745f646174615f62795f6c6f636b5f686173683137686361666239343538306137663634303645005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231345374616b65496e666f44656c7461313169735f696e6372656173653137683166386136356661303836623163316645005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231355374616b65417443656c6c446174613564656c74613137683762333332613765343438316530613845005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231345374616b65496e666f44656c746136616d6f756e743137683736303137613463316430633135626445005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231345374616b65496e666f44656c74613138696e61756775726174696f6e5f65706f63683137683538323561303933383837366165313345005f5a4e347574696c3668656c70657231376765745f63757272656e745f65706f63683137683561353332396138346166353437623445002e4c706372656c5f68693236002e4c706372656c5f68693237002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e3437002e4c706372656c5f68693234002e4c706372656c5f68693235002e4c616e6f6e2e63396664323635383763663061663763663065366537386464383734316533382e33002e4c706372656c5f68693239002e4c706372656c5f68693330002e4c706372656c5f68693331002e4c706372656c5f68693332002e4c706372656c5f68693333002e4c706372656c5f68693334002e4c706372656c5f68693335002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e34002e4c706372656c5f68693336007374722e30002e4c706372656c5f68693337007374722e31002e4c706372656c5f68693430002e4c706372656c5f68693339002e4c706372656c5f68693338005f5a4e34636f72653970616e69636b696e673970616e69635f666d74313768643661616165666234633464653863394500727573745f626567696e5f756e77696e64005f5a4e37636b625f7374643873797363616c6c73366e617469766534657869743137686334346330613764356530656238316345005f5a4e357374616b6531316f6f6d5f68616e646c65723137686231363437366264636564323636613345005f5f72675f6f6f6d005f5f72675f616c6c6f63005f5a4e3130365f244c542462756464795f616c6c6f632e2e6e6f6e5f746872656164736166655f616c6c6f632e2e4e6f6e54687265616473616665416c6c6f63247532302461732475323024636f72652e2e616c6c6f632e2e676c6f62616c2e2e476c6f62616c416c6c6f632447542435616c6c6f633137683966656332343337626566343266383945005f5f72675f6465616c6c6f63005f5a4e3130365f244c542462756464795f616c6c6f632e2e6e6f6e5f746872656164736166655f616c6c6f632e2e4e6f6e54687265616473616665416c6c6f63247532302461732475323024636f72652e2e616c6c6f632e2e676c6f62616c2e2e476c6f62616c416c6c6f6324475424376465616c6c6f633137686530336235656339643238613732396445005f5f72675f7265616c6c6f63005f5f72675f616c6c6f635f7a65726f6564005f5f727573745f616c6c6f63005f5f727573745f7265616c6c6f63005f5f727573745f616c6c6f635f7a65726f6564005f5f727573745f616c6c6f635f6572726f725f68616e646c6572005f5a4e35616c6c6f63377261775f766563313763617061636974795f6f766572666c6f773137683736396433373734353939336431626545002e4c706372656c5f68693431002e4c706372656c5f68693432002e4c706372656c5f68693433002e4c706372656c5f68693434002e4c706372656c5f68693435002e4c706372656c5f68693436002e4c706372656c5f68693437002e4c706372656c5f68693438005f5a4e396d6f6c6563756c65323672656164657238355f244c5424696d706c2475323024636f72652e2e636f6e766572742e2e46726f6d244c54246d6f6c6563756c65322e2e7265616465722e2e437572736f72244754242475323024666f7224753230247538244754243466726f6d3137686461653235633931336631613435396545002e4c706372656c5f68693439002e4c706372656c5f68693530002e4c706372656c5f68693531002e4c706372656c5f68693532005f5a4e396d6f6c6563756c65323672656164657238365f244c5424696d706c2475323024636f72652e2e636f6e766572742e2e46726f6d244c54246d6f6c6563756c65322e2e7265616465722e2e437572736f72244754242475323024666f722475323024753634244754243466726f6d3137686232663035653938653831303635333145002e4c706372656c5f68693533002e4c706372656c5f68693534002e4c706372656c5f68693535002e4c706372656c5f68693536002e4c706372656c5f68693537002e4c706372656c5f68693538005f5a4e3131626c616b6532625f7265663131626c616b6532625f7265663138626c616b6532625f696e69745f706172616d3137683431613831343963666239633164343445002e4c706372656c5f68693539005f5a4e3131626c616b6532625f7265663131626c616b6532625f7265663130626c616b6532625f49563137686532356438333932346363316638393145005f5a4e3131626c616b6532625f7265663131626c616b6532625f7265663134626c616b6532625f7570646174653137683337646637643338333264666265336545005f5a4e3131626c616b6532625f7265663131626c616b6532625f7265663136626c616b6532625f636f6d70726573733137683531363361326435303733336262323945002e4c43504932375f30002e4c43504932375f31002e4c43504932375f32002e4c43504932375f33002e4c43504932375f34002e4c43504932375f35002e4c43504932375f36002e4c43504932375f37002e4c706372656c5f68693630002e4c706372656c5f68693631002e4c706372656c5f68693632002e4c706372656c5f68693633002e4c706372656c5f68693634002e4c706372656c5f68693635002e4c706372656c5f68693636002e4c706372656c5f68693637005f5a4e313162756464795f616c6c6f63313162756464795f616c6c6f6331304275646479416c6c6f63336e65773137683039343964346234353436656265666245005f5a4e313162756464795f616c6c6f63313162756464795f616c6c6f6337726f756e6475703137686533656266373734346663663366363345002e4c706372656c5f68693735007374722e342e3336005f5a4e313162756464795f616c6c6f63313162756464795f616c6c6f63366e626c6f636b3137683537623963376462363561386133343745005f5a4e313162756464795f616c6c6f63313162756464795f616c6c6f6331304275646479416c6c6f633131626c6f636b5f696e6465783137683333633165376336333564613363643945005f5a4e34636f7265366f7074696f6e31336578706563745f6661696c65643137686332333330616533386638616564396545002e4c706372656c5f68693830002e4c706372656c5f68693736002e4c706372656c5f68693737002e4c706372656c5f68693638002e4c706372656c5f68693730007374722e322e3337002e4c706372656c5f68693731007374722e332e3338002e4c706372656c5f68693732002e4c706372656c5f68693733007374722e312e3335002e4c706372656c5f68693734002e4c706372656c5f68693831002e4c706372656c5f68693738007374722e302e3334002e4c706372656c5f68693639002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3135002e4c706372656c5f68693832002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3238005f5a4e34636f72653970616e69636b696e67313370616e69635f646973706c61793137683538303536323433613031393534316645002e4c706372656c5f68693739002e4c706372656c5f68693833002e4c706372656c5f68693834002e4c706372656c5f68693835002e4c706372656c5f68693836002e4c706372656c5f68693837002e4c706372656c5f68693839002e4c706372656c5f68693930002e4c706372656c5f68693838002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3338005f5a4e313162756464795f616c6c6f633130666173745f616c6c6f633946617374416c6c6f63336e65773137683239303962396561363461333531383845002e4c706372656c5f68693932002e4c706372656c5f68693931002e4c706372656c5f68693933002e4c706372656c5f68693934005f5a4e357374616b6535414c4c4f433137683937323962343239646165336531333345002e4c706372656c5f68693938002e4c706372656c5f6869313033002e4c706372656c5f6869313034002e4c706372656c5f6869313031002e4c706372656c5f6869313035002e4c706372656c5f6869313036002e4c706372656c5f6869313032002e4c706372656c5f68693937002e4c706372656c5f68693939002e4c706372656c5f6869313030002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e32002e4c706372656c5f68693935002e4c706372656c5f68693936002e4c706372656c5f6869313037002e4c706372656c5f6869313038002e4c706372656c5f6869313039002e4c706372656c5f6869313133002e4c706372656c5f6869313132002e4c706372656c5f6869313136002e4c706372656c5f6869313138002e4c706372656c5f6869313139002e4c706372656c5f6869313230002e4c706372656c5f6869313137002e4c706372656c5f6869313130002e4c706372656c5f6869313131002e4c706372656c5f6869313134002e4c706372656c5f6869313135005f5a4e35616c6c6f63377261775f7665633139526177566563244c54245424432441244754243131616c6c6f636174655f696e3137683334393639363464643031633234363645005f5a4e35616c6c6f63377261775f7665633139526177566563244c542454244324412447542437726573657276653231646f5f726573657276655f616e645f68616e646c653137686234636364626536643135363830353445002e4c706372656c5f6869313231007374722e302e3434005f5a4e35616c6c6f63377261775f7665633139526177566563244c5424542443244124475424313467726f775f616d6f7274697a65643137683131313435313531653037646531613245005f5a4e35616c6c6f63377261775f766563313166696e6973685f67726f773137683362363537323731663362336132663345005f5a4e35616c6c6f63377261775f7665633139526177566563244c54245424432441244754243136726573657276655f666f725f707573683137683364383734353931323332303230376445002e4c706372656c5f6869313232002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e313734002e4c706372656c5f6869313233002e4c706372656c5f6869313234005f5a4e36315f244c5424636b625f7374642e2e6572726f722e2e5379734572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137686534313062343262643137646531353845002e4c706372656c5f6869313235002e4c4a544934375f30002e4c424234375f31002e4c706372656c5f6869313236002e4c616e6f6e2e35366333623930656239393266643662383361623665306438306633656532622e3339002e4c424234375f32002e4c706372656c5f6869313237002e4c616e6f6e2e35366333623930656239393266643662383361623665306438306633656532622e3338002e4c424234375f33002e4c706372656c5f6869313238002e4c616e6f6e2e35366333623930656239393266643662383361623665306438306633656532622e3336002e4c706372656c5f6869313239002e4c616e6f6e2e35366333623930656239393266643662383361623665306438306633656532622e3337002e4c424234375f34002e4c706372656c5f6869313330002e4c424234375f36002e4c706372656c5f6869313331002e4c616e6f6e2e35366333623930656239393266643662383361623665306438306633656532622e3333002e4c706372656c5f6869313332002e4c616e6f6e2e35366333623930656239393266643662383361623665306438306633656532622e3334005f5a4e34636f726533666d7439466f726d6174746572323564656275675f7475706c655f6669656c64315f66696e6973683137683963326264643732306464613133376545005f5a4e34636f726533707472323864726f705f696e5f706c616365244c542424524624753634244754243137683135383466626334313265393865303445005f5a4e37636b625f7374643130686967685f6c6576656c31396c6f61645f63656c6c5f747970655f686173683137683563643636373336663632346636613545005f5a4e34636f7265336f70733866756e6374696f6e36466e4f6e63653963616c6c5f6f6e63653137683331326365396462383432326365623645005f5a4e34636f72653370747231303264726f705f696e5f706c616365244c542424524624636f72652e2e697465722e2e61646170746572732e2e636f706965642e2e436f70696564244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c542475382447542424475424244754243137683465633534623435323134663763393045002e4c43504935375f30005f5a4e34636f726533666d74336e756d33696d7037666d745f7536343137683238366534643532373433386334363745002e4c706372656c5f6869313333002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333234002e4c706372656c5f6869313334002e4c706372656c5f6869313335002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e3233005f5a4e34636f726533666d7439466f726d617474657231327061645f696e74656772616c3137686238656639343965396131613633346545005f5a4e34636f726533666d7439466f726d617474657231327061645f696e74656772616c313277726974655f7072656669783137683834663538656430383761336264393345002e4c43504936305f30002e4c43504936305f31005f5a4e34636f726533666d7439466f726d6174746572337061643137683433336537613934646232626438653245002e4c706372656c5f6869313336002e4c706372656c5f6869313337005f5a4e34636f726533666d743577726974653137683537653362636463656237646630393145002e4c706372656c5f6869313338005f5a4e36305f244c5424636f72652e2e63656c6c2e2e426f72726f774572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137686163386261333334363731373261333845002e4c706372656c5f6869313339002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e313730005f5a4e36335f244c5424636f72652e2e63656c6c2e2e426f72726f774d75744572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683636336332373865383138373636393045002e4c706372656c5f6869313430002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e313731005f5a4e34636f726533666d74336e756d35335f244c5424696d706c2475323024636f72652e2e666d742e2e4c6f7765724865782475323024666f7224753230246936342447542433666d743137686632356530653835343735353364373145002e4c706372656c5f6869313431002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333232002e4c43504936385f30002e4c43504936385f31002e4c43504936385f32005f5a4e36385f244c5424636f72652e2e666d742e2e6275696c646572732e2e50616441646170746572247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f7374723137686539366438303337316562386433343445002e4c706372656c5f6869313432002e4c706372656c5f6869313433002e4c706372656c5f6869313434002e4c706372656c5f6869313435005f5a4e34636f726533666d74355772697465313077726974655f636861723137686664666234386663643336373461323845005f5a4e34636f726533666d743557726974653977726974655f666d743137683364623431343565346436363932376245002e4c706372656c5f6869313436002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333237005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f7374723137683865303931326361326264646233386345005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e577269746524475424313077726974655f636861723137683239666437616639333939643762333645005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f666d743137683565373464633863623261616161323645002e4c706372656c5f6869313437005f5a4e34636f726533666d74386275696c64657273313044656275675475706c65356669656c643137686134393061356537663734366534656245002e4c706372656c5f6869313439002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e323933002e4c706372656c5f6869313530002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333030002e4c706372656c5f6869313438002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333031002e4c706372656c5f6869313531002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e323839002e4c706372656c5f6869313532002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e323932002e4c706372656c5f6869313534002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333032002e4c706372656c5f6869313533002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e313537005f5a4e34325f244c54242452462454247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137686332303631326561373836393861653445002e4c706372656c5f6869313535002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333337005f5a4e36375f244c5424636f72652e2e61727261792e2e54727946726f6d536c6963654572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683532646436363362353834636335356645002e4c706372656c5f6869313536002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e353537002e4c706372656c5f6869313537002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e353333002e4c706372656c5f6869313539002e4c706372656c5f6869313538005f5a4e34636f726533666d74336e756d35335f244c5424696d706c2475323024636f72652e2e666d742e2e55707065724865782475323024666f7224753230246936342447542433666d743137683464336136353331313038303933376445002e4c706372656c5f6869313630005f5a4e3133325f244c5424616c6c6f632e2e7665632e2e566563244c5424542443244124475424247532302461732475323024616c6c6f632e2e7665632e2e737065635f657874656e642e2e53706563457874656e64244c54242452462454244324636f72652e2e736c6963652e2e697465722e2e49746572244c5424542447542424475424244754243131737065635f657874656e643137683464663561353366366631653763336445005f5a4e35616c6c6f63377261775f7665633139526177566563244c542454244324412447542437726573657276653231646f5f726573657276655f616e645f68616e646c653137686332663335393562613638613033633645005f5a4e34325f244c54242452462454247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683431323134373832613466363464656645005f5a4e35616c6c6f63337665633136566563244c54245424432441244754243131657874656e645f776974683137683935323361376565386561616133316645005f5a4e35616c6c6f63377261775f7665633139526177566563244c542454244324412447542437726573657276653231646f5f726573657276655f616e645f68616e646c653137686534386235666233366361343936633545005f5a4e35616c6c6f63377261775f766563313166696e6973685f67726f773137686465323762646133633136313431313345005f5a4e396d6f6c6563756c65323672656164657237726561645f61743137686436323832346538376630396538383045002e4c706372656c5f6869313730007374722e312e323739002e4c706372656c5f6869313633002e4c706372656c5f6869313634002e4c706372656c5f6869313631002e4c706372656c5f6869313632002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e31002e4c706372656c5f6869313639002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3136002e4c706372656c5f6869313731002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3139002e4c706372656c5f6869313635002e4c706372656c5f6869313636002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e36002e4c706372656c5f6869313637002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3132002e4c706372656c5f6869313638002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3134005f5a4e36315f244c54246d6f6c6563756c65322e2e7265616465722e2e4572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683238346238363235356264316239336545002e4c706372656c5f6869313732002e4c7377697463682e7461626c652e5f5a4e36315f244c54246d6f6c6563756c65322e2e7265616465722e2e4572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683238346238363235356264316239336545002e4c706372656c5f6869313733002e4c7377697463682e7461626c652e5f5a4e36315f244c54246d6f6c6563756c65322e2e7265616465722e2e4572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d7431376832383462383632353562643162393365452e333539005f5a4e396d6f6c6563756c65323672656164657236437572736f723876616c69646174653137683930306131623931383065653939313845002e4c706372656c5f6869313736002e4c706372656c5f6869313734002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e32002e4c706372656c5f6869313735002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e33002e4c706372656c5f6869313737002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3238005f5a4e396d6f6c6563756c65323672656164657236437572736f723133756e7061636b5f6e756d6265723137683635326430373132666263326536343145002e4c706372656c5f6869313738002e4c706372656c5f6869313739002e4c706372656c5f6869313830002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3331002e4c706372656c5f6869313831002e4c706372656c5f6869313839002e4c706372656c5f6869313832002e4c706372656c5f6869313833002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3335002e4c706372656c5f6869313834002e4c706372656c5f6869313838002e4c706372656c5f6869313835002e4c706372656c5f6869313836002e4c706372656c5f6869313837002e4c706372656c5f6869313930002e4c706372656c5f6869313931002e4c706372656c5f6869313932002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3430002e4c706372656c5f6869313933002e4c706372656c5f6869313934002e4c706372656c5f6869313935002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3538002e4c706372656c5f6869313936002e4c706372656c5f6869313937002e4c706372656c5f6869313938002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3634005f5a4e36395f244c5424616c6c6f632e2e7665632e2e566563244c54247538244754242475323024617324753230246d6f6c6563756c65322e2e7265616465722e2e526561642447542434726561643137683538323363346134366134643066373445002e4c706372656c5f6869313939002e4c706372656c5f6869323030002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3638005f5a4e34636f726533707472343664726f705f696e5f706c616365244c5424616c6c6f632e2e7665632e2e566563244c5424753824475424244754243137683139303635656264313265376238616645002e4c706372656c5f6869323031005f5a4e3130325f244c5424636f72652e2e697465722e2e61646170746572732e2e6d61702e2e4d6170244c5424492443244624475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424387472795f666f6c643137686639333339613334663266393033663145002e4c706372656c5f6869323035002e4c706372656c5f6869323034002e4c706372656c5f6869323032002e4c706372656c5f6869323033002e4c706372656c5f6869323036002e4c4a54493130335f30002e4c42423130335f31002e4c42423130335f32002e4c42423130335f33002e4c42423130335f34002e4c42423130335f35002e4c706372656c5f6869323134002e4c706372656c5f6869323039007374722e322e3433002e4c706372656c5f6869323130002e4c706372656c5f6869323131002e4c706372656c5f6869323132002e4c706372656c5f6869323133002e4c706372656c5f6869323037002e4c706372656c5f6869323038002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e3439002e4c706372656c5f6869323136002e4c706372656c5f6869323135002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e313133002e4c706372656c5f6869323137002e4c706372656c5f6869323138002e4c706372656c5f6869323139002e4c706372656c5f6869323230002e4c706372656c5f6869323231002e4c706372656c5f6869323232002e4c616e6f6e2e62303761633263373733636532303537336637343863366132643634626130332e313138002e4c706372656c5f6869323233005f5a4e357374616b6531315f42554444595f484541503137683738323931303732643365343635303345005f5a4e357374616b6531375f46495845445f424c4f434b5f484541503137686366636131376364336532396638393845002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3134002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3237002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3732002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3733002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3734002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3735002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3736002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3737002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3738002e4c6c696e655f7461626c655f737461727430002e4c6c696e655f7461626c655f737461727431006c69622e63002478002478002478002478002e4c32002e4c33002e4c3335002e4c3437002e4c3132002e4c3739002e4c3830002e4c3134002e4c3135002e4c3136002e4c3831002e4c3138002e4c3230002e4c3231002e4c3738002e4c3235002e4c3236002e4c3237002e4c3238002e4c3331002e4c3332002e4c3333002e4c3334002e4c3330002e4c3137002e4c3239002e4c3130002e4c313433002e4c313437002e4c313438002e4c313439002e4c323033002e4c313532002e4c323034002e4c313735002e4c313736002e4c313632002e4c323031002e4c313737002e4c313638002e4c313730002e4c313738002e4c313731002e4c313733002e4c313536002e4c313539002e4c313630002e4c313631002e4c313634002e4c323035002e4c313537002e4c313637002e4c313534005f5f636b625f7374645f6d61696e005f7374617274006d656d736574006d656d637079006d656d636d70006d656d6d6f7665000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000120000000000000060010100000000006001000000000000680900000000000000000000000000001000000000000000000000000000000009000000010000000200000000000000c80a010000000000c80a0000000000001c0c00000000000000000000000000000800000000000000000000000000000013000000010000000600000000000000e426010000000000e416000000000000fa8400000000000000000000000000000400000000000000000000000000000019000000010000000300000000000000e0bb010000000000e09b00000000000070000000000000000000000000000000080000000000000000000000000000002000000001000000030000000000000050bc010000000000509c000000000000b8000000000000000000000000000000080000000000000000000000000000002600000008000000030000000000000008bd010000000000089d00000000000000200800000000000000000000000000010000000000000000000000000000002b0000000100000000000000000000000000000000000000089d0000000000000c02000000000000000000000000000001000000000000000000000000000000390000000100000000000000000000000000000000000000149f0000000000001b230000000000000000000000000000010000000000000000000000000000004500000001000000000000000000000000000000000000002fc2000000000000f0010000000000000000000000000000010000000000000000000000000000005400000001000000000000000000000000000000000000001fc400000000000020100000000000000000000000000000010000000000000000000000000000006200000001000000300000000000000000000000000000003fd4000000000000274c0000000000000000000000000000010000000000000001000000000000006d00000001000000000000000000000000000000000000006620010000000000171b0000000000000000000000000000010000000000000000000000000000007d00000001000000000000000000000000000000000000007d3b01000000000024000000000000000000000000000000010000000000000000000000000000008d0000000300007000000000000000000000000000000000a13b0100000000002b000000000000000000000000000000010000000000000000000000000000009f0000000100000000000000000000000000000000000000cc3b0100000000004c1c000000000000000000000000000001000000000000000000000000000000ab000000010000003000000000000000000000000000000018580100000000002300000000000000000000000000000001000000000000000100000000000000b40000000200000000000000000000000000000000000000405801000000000050e2000000000000130000006c09000008000000000000001800000000000000bc0000000300000000000000000000000000000000000000903a020000000000ce00000000000000000000000000000001000000000000000000000000000000c600000003000000000000000000000000000000000000005e3b0200000000001d3a000000000000000000000000000001000000000000000000000000000000",
        "0x"
      ],
      "witnesses": [
        "0x5500000010000000550000005500000041000000be5098c531d52a249e691b627e5eea2d195178f2072eeda1d4c7b4d87fd018bd310b83981d8bb6da7e5c5110040da5c1eac2b480ac12f88eb83228d5c99004d801"
      ]
    }
  },
  "cell_tx": {
    "version": "0x0",
    "cell_deps": [
      {
        "out_point": {
          "tx_hash": "0xf8de3bb47d055cdf460d93a2a6e1b05f7432f9777c8c474abf4eec1d4aee5d37",
          "index": "0x0"
        },
        "dep_type": "dep_group"
      }
    ],
    "header_deps": [],
    "inputs": [
      {
        "since": "0x0",
        "previous_output": {
          "tx_hash": "0xbe3777fa551ec2de85ece9cca9918eefc953db190d52426d74c5f1cc73b2868c",
          "index": "0x1"
        }
      },
      {
        "since": "0x0",
        "previous_output": {
          "tx_hash": "0xe6a4b80a06bbfbdb23456e6845b8ee87aa9644ad185c25295c919dbe6dbd8da0",
          "index": "0x1"
        }
      }
    ],
    "outputs": [
      {
        "capacity": "0xed2b86be600",
        "lock": {
          "code_hash": "0x9bd7e06f3ecf4be0f2fcd2188b23f1b9fcc88e5d4b65a8637b17723bbda3cce8",
          "hash_type": "type",
          "args": "0x61a0d1fa2b4a4536a778659d5d87b88e82188b17"
        },
        "type": {
          "code_hash": "0x00000000000000000000000000000000000000000000000000545950455f4944",
          "hash_type": "type",
          "args": "0xb7fe83392736c6d1633f35194d1a0e7e87fcc908a84394074031b5b95e06c026"
        }
      },
      {
        "capacity": "0x18591bf1fe00",
        "lock": {
          "code_hash": "0x9bd7e06f3ecf4be0f2fcd2188b23f1b9fcc88e5d4b65a8637b17723bbda3cce8",
          "hash_type": "type",
          "args": "0x61a0d1fa2b4a4536a778659d5d87b88e82188b17"
        },
        "type": {
          "code_hash": "0x00000000000000000000000000000000000000000000000000545950455f4944",
          "hash_type": "type",
          "args": "0xf89735de346f9655e16d60c3d91963fe67f8b845f511e5fcdea60d462c94a33e"
        }
      },
      {
        "capacity": "0x12d9e4a31c3fd",
        "lock": {
          "code_hash": "0x9bd7e06f3ecf4be0f2fcd2188b23f1b9fcc88e5d4b65a8637b17723bbda3cce8",
          "hash_type": "type",
          "args": "0x61a0d1fa2b4a4536a778659d5d87b88e82188b17"
        },
        "type": null
      }
    ],
    "outputs_data": [
      "0x7f454c460201010000000000000000000200f30001000000d426010000000000400000000000000028770200000000000100000040003800050040001400120006000000040000004000000000000000400001000000000040000100000000001801000000000000180100000000000008000000000000000100000004000000000000000000000000000100000000000000010000000000d416000000000000d41600000000000000100000000000000100000005000000d416000000000000d426010000000000d4260100000000001c850000000000001c8500000000000000100000000000000100000006000000f09b000000000000f0bb010000000000f0bb01000000000028010000000000002821080000000000001000000000000051e574640600000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c740100000000005e74010000000000707401000000000088740100000000009e7401000000000020950100000000001e95010000000000229501000000000026950100000000002a95010000000000c874010000000000000000000000000001000000000000003686010000000000617474656d707420746f206164642077697468206f766572666c6f7700000000617474656d707420746f2073756274726163742077697468206f766572666c6f7700000000000000c87401000000000001000000000000000100000000000000088c01000000000008c9bcf367e6096a3ba7ca8485ae67bb2bf894fe72f36e3cf1361d5f3af54fa5d182e6ad7f520e511f6c3e2b8c68059b6bbd41fbabd9831f79217e1319cde05bc874010000000000000000000000000001000000000000000c800100000000000000000000000000617474656d707420746f207368696674206c6566742077697468206f766572666c6f7700000000000000000000000000617474656d707420746f206d756c7469706c792077697468206f766572666c6f77000000000000000000000000000000617474656d707420746f2073756274726163742077697468206f766572666c6f77000000000000000000000000000000617474656d707420746f2073686966742072696768742077697468206f766572666c6f77000000000000000000000000617474656d707420746f206164642077697468206f766572666c6f776c6561662073697a65206d75737420626520616c69676e20746f203136206279746573007c0301000000000023000000000000007265717569726573206d6f7265206d656d6f727920737061636520746f20696e697469616c697a65204275646479416c6c6f630000000000b00301000000000033000000000000006f7574206f66206d656d6f72790000000000000000000000617474656d707420746f20646976696465206279207a65726f00000000000000617474656d707420746f206164642077697468206f766572666c6f77427974655265616465724279746533325265616465724279746573526561646572000000617474656d707420746f2073756274726163742077697468206f766572666c6f775363726970745265616465725769746e65737341726773526561646572556e6b6e6f776e000000c874010000000000080000000000000008000000000000007a88010000000000456e636f64696e674f766572666c6f7776616c69646174654c656e6774684e6f74456e6f75676800c874010000000000080000000000000008000000000000007a880100000000004974656d4d697373696e67496e6465784f75744f66426f756e6429426f72726f774572726f72426f72726f774d75744572726f7200000000787701000000000018000000000000000800000000000000b880010000000000748201000000000028830100000000002020202052656164446174612c0a2c20280a282c30783030303130323033303430353036303730383039313031313132313331343135313631373138313932303231323232333234323532363237323832393330333133323333333433353336333733383339343034313432343334343435343634373438343935303531353235333534353535363537353835393630363136323633363436353636363736383639373037313732373337343735373637373738373938303831383238333834383538363837383838393930393139323933393439353936393739383939000078770100000000000800000000000000080000000000000060830100000000006a8301000000000020840100000000002829000000000000787701000000000008000000000000000800000000000000208601000000000054727946726f6d536c6963654572726f72636b622d64656661756c742d68617368616c726561647920626f72726f77656400000000000000c874010000000000000000000000000001000000000000000c80010000000000616c7265616479206d757461626c7920626f72726f776564c87401000000000000000000000000000100000000000000fa7f01000000000063616c6c656420604f7074696f6e3a3a756e77726170282960206f6e206120604e6f6e65602076616c75650000000000c87401000000000001000000000000000100000000000000088c010000000000617474656d707420746f206164642077697468206f766572666c6f77726561645f6174206069662073697a65203c20726561645f6c656e60726561645f6174206069662064732e63616368655f73697a65203e2064732e6d61785f63616368655f73697a6560726561645f617420606966206375722e6f6666736574203c2064732e73746172745f706f696e74207c7c202e2e2e60726561645f61742060696620726561645f706f696e74202b20726561645f6c656e203e2064732e63616368655f73697a656076616c69646174653a2073697a65203e206375722e736f757263652e746f74616c5f73697a65756e7061636b5f6e756d6265726765745f6974656d5f636f756e74636f6e766572745f746f5f753634636f6e766572745f746f5f7538636f6e7665727420746f205665633c75383e00000096910100000000001800000000000000080000000000000062900100000000004669656c64436f756e744f75744f66426f756e64556e6b6e6f776e4974656d4f6666736574486561646572546f74616c53697a65436f6d6d6f6e0000000000000000000000000000617474656d707420746f206164642077697468206f766572666c6f770000000063616c6c65642060526573756c743a3a756e77726170282960206f6e20616e2060457272602076616c75650000000000c874010000000000000000000000000001000000000000003686010000000000c874010000000000100000000000000008000000000000003674010000000000617373657274696f6e206661696c65643a20636865636b706f696e745f646174612e69735f6e6f6e652829617373657274696f6e206661696c65643a207374616b655f61745f646174612e69735f6e6f6e6528290000000006000000000000000900000000000000060000000000000006000000000000000b000000000000000a000000000000000a000000000000000400000000000000080000000000000004000000000000002c0901000000000023090100000000001d0901000000000017090100000000000c090100000000000209010000000000f8080100000000009005010000000000e0040100000000008c050100000000001000000000000000017a5200017801011b0c02002c00000018000000061c0000181b000000440ed00d74810188028903920493059406950796089709980a990b9a0c9b0d1000000048000000ee3600000a000000000e0000100000005c000000e436000008000000000000001000000070000000d836000008000000000000001c00000084000000cc3600004e00000000420e304a810188028903920493050018000000a4000000fa3600003000000000420e20468101880289030014000000c00000000e3700000e00000000420e104281010014000000d8000000043700000e00000000420e104281010018000000f0000000fa3600005800000000420e404481018802000000180000000c010000363700005800000000420e4044810188020000001800000028010000723700005800000000420e4044810188020000001800000044010000ae3700005800000000420e4044810188020000001400000060010000ea3700005200000000420e40428101001800000078010000243800005800000000420e4044810188020000001400000094010000603800005200000000420e404281010018000000ac0100009a3800005800000000420e40448101880200000018000000c8010000d63800004e00000000420e3044810188020000001c000000e4010000083900009a00000000420e20488101880289039204000000200000000402000082390000dc00000000440e304c8101880289039204930594060000002c000000280200003a3a0000ee1a000000420ef0035a810188028903920493059406950796089709980a990b9a0c9b0d2c00000058020000f85400001404000000420e80015a810188028903920493059406950796089709980a990b9a0c9b0d1000000088020000dc5800003c000000000e0000100000009c020000045900000a000000000e000010000000b0020000fa5800004c000000000e000010000000c4020000325900004c000000000e000010000000d80200006a590000f4000000000e00002c000000ec0200004a5a0000d403000000420eb00158810188028903920493059406950796089709980a990b9a0c00002c0000001c030000ee5d0000f203000000420ec0015a810188028903920493059406950796089709980a990b9a0c9b0d200000004c030000b0610000d600000000420e504e8101880289039204930594069507001800000070030000626200005200000000420e204681018802890300140000008c030000986200003400000000420e104281010018000000a4030000b46200007400000000420e50468101880289030014000000c00300000c6300003600000000420e104281010020000000d80300002a6300006c00000000420e304c81018802890392049305940600000020000000fc030000726300006200000000420e304c8101880289039204930594060000001000000020040000b063000022000000000e00001800000034040000be6300003a00000000420e2046810188028903002000000050040000dc630000fc00000000420e404e8101880289039204930594069507001000000074040000b464000042000000000e00001400000088040000e26400009200000000420e104281010010000000a00400005c650000020000000000000010000000b40400004a650000360000000000000018000000c80400006c6500007a00000000420e40448101880200000018000000e4040000ca6500008200000000420e4044810188020000002400000000050000306600006001000000440ee0086481018802890392049305940695079608970910000000280500006867000018000000000e0000100000003c0500006c670000040000000000000010000000500500005c670000020000000000000014000000640500004a6700004201000000420e30428101002c0000007c05000074680000e401000000420e705a810188028903920493059406950796089709980a990b9a0c9b0d001c000000ac050000286a00005600000000420e304a810188028903920493050024000000cc0500005e6a00007803000000420e50528101880289039204930594069507960897090014000000f4050000ae6d00000e00000000420e1042810100240000000c060000a46d00007e01000000420e8001508101880289039204930594069507960800001000000034060000fa6e000012000000000000001000000048060000f86e00001200000000000000140000005c060000f66e00000e00000000420e10428101001400000074060000ec6e00000e00000000420e1042810100140000008c060000e26e00000e00000000420e104281010014000000a4060000d86e00007000000000420e90014281012c000000bc060000306f0000bc01000000420e90015a810188028903920493059406950796089709980a990b9a0c9b0d14000000ec060000bc700000b400000000420e10428101001400000004070000587100003800000000420e4042810100100000001c070000787100000a0000000000000014000000300700006e710000b600000000420e104281010014000000480700000c7200003a00000000420e404281010020000000600700002e7200002001000000420ea0014e81018802890392049305940695071c000000840700002a7300009800000000420e4048810188028903920400000014000000a4070000a27300000e00000000420e104281010010000000bc07000098730000160000000000000018000000d00700009a730000a200000000420e40468101880289030014000000ec070000207400007000000000420e90014281011c00000004080000787400005200000000420e304a81018802890392049305001800000024080000aa7400007e00000000420e5046810188028903001c000000400800000c7500006200000000420e2048810188028903920400000010000000600800004e750000300000000000000018000000740800006a7500004e00000000420e1044810188020000001c000000900800009c7500006800000000420e304a810188028903920493050018000000b0080000e47500007e00000000420e50468101880289030018000000cc080000467600005200000000420e20468101880289030018000000e80800007c7600005600000000420e1044810188020000002000000004090000b67600008201000000420e504e8101880289039204930594069507001000000028090000147800002800000000000000100000003c090000287800006200000000420e101800000050090000767800006800000000420e304481018802000000180000006c090000c27800005400000000420e3044810188020000002400000088090000fa7800007c01000000420e80015281018802890392049305940695079608970918000000b00900004e7a00007800000000420e40468101880289030018000000cc090000aa7a00007e00000000420e4046810188028903001c000000e80900000c7b0000a200000000420e5048810188028903920400000018000000080a00008e7b00007a00000000420e20468101880289030020000000240a0000ec7b0000ba00000000420e504c81018802890392049305940600000010000000480a0000827c00001000000000000000100000005c0a00007e7c0000080000000000000010000000700a0000727c0000080000000000000010000000840a0000667c0000080000000000000010000000980a00005a7c0000080000000000000010000000ac0a00004e7c00000a000000000e00001c000000c00a0000447c00007200000000420e5048810188028903920400000024000000e00a0000967c0000ca02000000420ea0015081018802890392049305940695079608000010000000080b0000387f000028000000000e0000240000001c0b00004c7f00006401000000420ea0015081018802890392049305940695079608000024000000440b0000888000008605000000440e800864810188028903920493059406950796089709280000006c0b0000e68500001803000000420eb00256810188028903920493059406950796089709980a990b18000000980b0000d28800009200000000420eb001468101880289032c000000b40b000048890000a003000000420ed0025a810188028903920493059406950796089709980a990b9a0c9b0d24000000e40b0000b88c00008601000000420e90014c8101880289039204930594060000000000000000000002452c00014697000000e78000019308d00573000000130101932334116c2330816c233c916a2338216b2334316b2330416b233c5169233861692334716923308169233c91672338a1672334b167179600001306665e0ce208e6080c1306004013040040814597800000e78040db2338816205659b08458093050163080c09440146814601478147014873000000aa84630285080545638da406114463900418033b01631305004063786507854505445a8597600000e7804012aa8cae8a0c0c1306004097800000e78040e293020bc013850c402338516285659b88458093050163130600400943814601478147014873000000630d6510aa846309851011446397041083340163094463e29210a1a0014429a2054419a25a85814597600000e780a00baa8cae8a0c0c5a8697800000e780c0db114463708b023145b14b814597600000e78060092a892e8a17e5ffff930515c791a003c51c0083c50c0003c62c0083c63c0022054d8d4206e206558e3364a600631a8b02214463788b0e3145b14b814597600000e78020052a892e8a17e5ffff9305d5c231464a8597800000e780c0d485442da03145b14b814597600000e78080022a892e8a17e5ffff930535c031464a8597800000e78020d28144da8923289120232a8121233c8120233031232334212323384123233c7123080c97500000e78060c00d4463870a00668597700000e780a08dda8409a8014463870a00668597700000e780608c2285a68597700000e78080c12a841315840361958330816c0334016c8334816b0339016b8339816a033a016a833a8169033b0169833b8168033c0168833c8167033d0167833d81661301016d828003c55c0083c54c0003c66c0083c67c0022054d8d4206e206558e3364a6001335840093753400b335b0004d8d15c531453149814597600000e78080f32a84ae8917e5ffff930535b13146228597800000e78020c38d4409bf63708b023145b14b814597600000e780a0f02a892e8a17e5ffff930555ae65bd93592400fd190d4563f8a9023145b14b814597600000e78020ee2a892e8a17e5ffff9305d5ab31464a8597800000e780c0bd91440d446dbd639ea908114691446685da85a28697500000e780008a13f63500f199b306b5002338a120233cb1202330d1222334c12223389122130501630c0c97400000e780005a13050163da8597500000e7808088033901638334016423382121233c912009452330a122080c97500000e780e09921cd31453149814597600000e78040e42a84ae8917e5ffff9305f5a13146228597800000e780e0b38d4459aa3145b14b814597600000e780a0e12a892e8a17e5ffff9305559f31464a8597800000e78040b10d449144cdbb6380047605456380a47603360900833689006685da8597400000e780007d13040002639e850e09456382a47403368900833609016685da8597400000e780e07a0544639e850e0d456385a47203360901833689016685da8597400000e780e0782a86ae86080cb285368697400000e780807d8324012115456393a4100335816311c54a8597600000e78040672d45636465016f10e00d93054bff0d456364b5006f10c00403c5dc0083c5cc0003c6ec0083c6fc0022054d8d4206e206558e83c51c0083c60c0003c72c0083873c00a205d58d4207e2075d8fd98d1147b366a600638ce50a03c55c0083c54c0003c66c0003877c0022054d8d42066207598e518d8d4563f6a56a7199c1456317b508080ce6855a8697400000e78000674da8ae893145b14b814597600000e780e0cc2a892e8a17e5ffff9305e586314605a0ae892945a94b814597600000e780e0ca2a892e8a17e5ffff9305458429464a8597800000e780809a814403358163e30205c80335016397600000e780405895b9032c4121033481218339012203398122033a0123833b8123c9bf93050bff0d45e377b57403c51c0183c50c0103c62c0103c73c0122054d8d42066207598e3367a600080ce6855a8697400000e78020550334012103360122281a9146a28597400000e780805a0335812111c5228597600000e780c0507279b6642685814597600000e78080bf2a84ae89ca85268697800000e780a08f23388120233c312123309122130501630c0c97600000e780004003390163033481631305016313070002ca852286814697600000e780000003350163e30405720335016483358163033601632330a122233cb1202338c120880a0c0c97600000e780a02913050163930600025147ca85228697600000e780e0fb03350163e30c056e0335016483358163033601632330a122233cb1202338c120a8120c0c97600000e7808025080c1306004013040040814597700000e78020772338816205659b08a581054562151307150093050163080c01468146814701487300000021c54944567511c5367597600000e780c03f766511c5566597600000e780e03e4a8597600000e78060c6166511c5727597600000e780603de38f0ab0668597600000e780803c01be033a0163130510406367aa0685450544528597600000e78080aaaa892efa0c0c1306004097700000e780807a93040ac0138509402338916285659b88a581131784030507930501631306004081468147014873000000833501633335a000b3b5b4004d8d21c9527529d94e8597600000e780203599b75285814597600000e78000a4aa892efa0c0c528697700000e7802074114463708a024545454c814597600000e780c0a12a8bae8b17d5ffff9305356091a003c5190083c5090003c6290083c6390022054d8d4206e206558e3364a600631a8a02214463788a084545454c814597600000e780809d2a8bae8b17d5ffff9305f55b45465a8597700000e780206d054d2da04545454c814597600000e780e09a2a8bae8b17d5ffff9305555945465a8597700000e780806a014d2328a121232ab121233c8120233041232334612323387123233c8123080c97400000e780e05849445275e30205e64e8597600000e780002699bd03c5590083c5490003c6690083c6790022054d8d4206e206558e3364a6001335840093753400b335b0004d8d15c54545454b814597600000e780e0912a842e8a17d5ffff930555504546228597700000e78080610d4d85bf63708a024545454c814597600000e780008f2a8bae8b17d5ffff9305754d21bf93542400fd140d4563f8a4024545454c814597600000e780808c2a8bae8b17d5ffff9305f54a45465a8597700000e780205c114d0d44e1a0639ea408114691444e85d285a28697400000e780602813f63500f199b306b5002338a120233cb1202330d1222334c12223389122130501630c0c97400000e78060f813050163d28597400000e780e026033b01630334016423386121233c812009452330a122080c97400000e780403829cd4545454b814597600000e780a0822a842e8a17d5ffff930515414546228597700000e78040520d4d75a24545454c814597600000e78000802a8bae8b17d5ffff9305753e45465a8597700000e780a04f0d44114d268ab9b56302041405456302a41403360b0083368b004e85d28597400000e780401b99cd2a86ae86080cb285368697400000e780c01f032d012115456316ad1209456309a41003368b0083360b014e85d28597400000e780c01799cd2a86ae86080cb285368697400000e780401c032d01211545631aad0e0d456300a40e03360b0183368b014e85d28597400000e780401499cd2a86ae86080cb285368697400000e780c018032d01211545631ead0a0335816311c55a8597600000e780800293058aff0d45e377b52093054affe373b52003c5990083c5890003c6a90083c6b90022054d8d4206e206558eb366a60003c5d90083c5c90003c6e90003c7f90022054d8d42066207598e3367a600080cce85528697400000e780c0fe033501222aee49c503340121f2642685814597500000e780e06a2a8a2eeaa285268697700000e780003ba5a00145814509a80545854531a00945894519a00d458d4597500000e780603e0000832d412103348121033a0122033b8122833b0123033c812303358163e30605cc0335016397600000e78040f575b917d5ffff1305c5209305100297500000e780e0bf0000014a0335812119c50335012197600000e78080f263080a3a0d45f265e37cb55a03451a0083450a0003462a0083063a0022054d8d4206e206558e518d854529446318b554167593050002e31fb568d667014b02f603c5970183c5870103c6a70183c6b70122054d8d4206e206558e518d83c5d70103c6c70183c6e70103c7f701a205d18dc2066207d98ed58d82154d8daae303c5170183c5070103c6270183c6370122054d8d4206e206558e518d83c5570103c6470183c6670103c77701a205d18dc2066207d98ed58d82154d8d2aff03c5970083c5870003c6a70083c6b70022054d8d4206e206558e518d83c5d70003c6c70083c6e70003c7f700a205d18dc2066207d98ed58d82154d8d2afb03c5170083c5070003c6270083c6370022054d8d4206e206558e518d83c5570003c6470083c667003ee603c77700a205d18dc2066207d98ed58d82154d8d2af70d45aaff23300120130d1121930d9165080cac1b97600000e78040df034501218945630cb5246303051003459d0183458d010346ad018346bd0122054d8d4206e206558e518d8345dd010346cd018346ed010347fd01a205d18dc2066207d98ed58d82154d8d2334a16403451d0183450d0103462d0183463d0122054d8d4206e206558e518d83455d0103464d0183466d0103477d01a205d18dc2066207d98ed58d82154d8d2330a16403459d0083458d000346ad008346bd0022054d8d4206e206558e518d8345dd000346cd008346ed000347fd00a205d18dc2066207d98ed58d82154d8d233ca16203451d0083450d0003462d0083463d0022054d8d4206e206558e518d83455d0003464d0083466d0003477d00a205d18dc2066207d98ed58d82154d8d2338a16209a82334016423300164233c016223380162130501632c131306000297700000e780604d012519c1b27419aa130501630d46da8597400000e780600d03340163e301042e033581632af2833401642685814597500000e7806036aa8b2e8ca285268697700000e780800623387163233c816323309164130501659305016397600000e780c0b60385ed008385dd0003c6cd0083340165230fa162a205d18d231eb16203c59d0083c58d0003c6ad008386bd0022054d8d4206e206558e518d232ca16203c51d0083c50d0003c62d0083c63d0022054d8d4206e20683c55d00558e518d03c64d00a20583c66d0003c77d00d18d834b8165c2066207d98ed58d82154d8d2338a162327511c5327597500000e78020430305e1638315c16303268163833601632307a11e2316b11e2324c11eb6f3127511c5228597600000e78040b87d556300ab56050b26f671bb294419b232756301051c0305e11e8315c11e0326811e9e76230ba11c231ab11c2328c11cb6e713051162ac033d4697700000e78000f53275233ca16023007163080c930581610d4697500000e780806c033b0121e3010b2e0305712283056122034651222303a11aa205d18d2312b11a0345212283451122034631228306412222054d8d4206e206558e518d2320a11a0345a121834591210346b1218346c12122054d8d4206e2068345e121558e518d0346d121a2058346f12103470122d18d03048121c2066207d98ed58d82154d8d2aef327597500000e780e031130591182c0b3d4697700000e780a0e95ae323048118130501630c030d4697500000e780606103350163e30505240335016483358163033601632330a122233cb1202338c12028130c0c97600000e780c085130501630c03114697500000e780a05d03350163e30005220335016483358163033601632330a122233cb1202338c120130501630c0c97600000e780e081ba7d7a768334016303370164080cee85a68697600000e780c0ed0c0c13060002326597700000e7808021833581632a8491c5268597600000e780009d5a7511c56e8597600000e780209c0dc45a8597500000e78080231304300319a01304b0065265630d05f2528597600000e780c0996ff0cff2080c9146d285726697400000e78040a1833b0121833401222685814597500000e78000072a842e8bde85268697700000e78020d7e38004168344040063070b00228597600000e780e0940335812119c50335012197600000e780c093526511c5528597600000e780e0920545638aa4024944639b042e080c0546814597400000e78060c60345012163090510033581218335012297600000e780a0c52a84e9a4130501650c0397100000e780a0af28130c0397100000e780e0a3130501630c0397100000e78080a83a747a768334016303370164080ca285a68697600000e78000da13050002814597500000e78040faaa8b2e8b0c0c1306000297700000e78040ca0335816311c5268597600000e78060885a7511c5228597600000e780808793050002054685445e8597700000e78000a21375f50f13043004631e95029305000209465e8597700000e78040a01375f50f13044004631095028334016583350166268597600000e78020bb2a841375f50f630c052063070b005e8597600000e7804081033581656300051e0335016597600000e7800080c1aa0305712183056121034651212307a11aa205d18d2316b11a0345212183451121034631218306412122054d8d4206e206558e518d2324a11a033581228305012303348121833401222338a162230cb1621305f11b93050163254697700000e780a0ba13558403230ba11a13550403a30aa11a13558402230aa11a13550402a309a11a135584012309a11a13550401a308a11a135584002308a11aa307811a13d58403230fa11a13d50403a30ea11a13d58402230ea11a13d50402a30da11a13d58401230da11a13d50401a30ca11a13d58400230ca11aa30b911a130501650c0397100000e780a0a7080c0c0397100000e78020810334016503360166833401210337012213050163a285a68697600000e78040bd0335812111c5268597500000e780a06d0335816511c5228597500000e780a06c13050002814597500000e78080dbaa8d2e8b930501631306000297700000e78060aba8030c0397100000e780c08a3e65fe6597600000e78060a12a841375f50f05ed080cac03054697600000e78020400345012105e10334812283340122080cac03094697600000e780603e0345012163020510034411215e6511c53e6597500000e780406463070b006e8597500000e78060631375f40f29c11a6597500000e78080ea6ff06fbb17d5ffff1305c5daf1456ff02fed11456ff08fe863070b005e8597500000e78000600335816511c5268597500000e780005f1a6597500000e78080e6527511c54e8597500000e780805d567511c5367597500000e780a05c766511c5566597500000e780c05b4a8597500000e78040e3166511c5727597500000e780405a63870a00668597500000e780605901446fe0dfcd3145da856ff02fe017d5ffff130525d397c5ffff9386255e09a817d5ffff130505d297c5ffff9386055d9305b002100c97400000e780803c00000335012283358122258da18d4d8d3d44e31a05ee080c2c13054697600000e780e034833b012263880b0c033581212af60335812283350123033681238336012136f22338a164233cb1642330c166aefbaaf7def3080c2c13094697600000e780e030033c0122630b0c08033581212aee0335812283350123033681238336012136ea2338a164233cb1642330c1662334b1202330a120e2ff881397000000e780c0719374f50fa81b97000000e780e0701375f50f51446399a43c130501658c1397000000e780207f080cac1b97000000e780607e03360166033501226313a602833501210335016597700000e780c0c9133a150001a80344012129b50344012149ae014a0335812119c50335012197500000e78000440335816519c50335016597500000e780e04263000a36130581618c1397000000e780807d080c9305816197000000e780806c8335012241456397a54403350121834585002ee583459500aefc8345a500aef88345b500aef48345c500aef08345d5002efc8345e5002ef88345f5002ef4834505002ee183451500aeec83452500aee883453500aee483454500aee0834555002ef0834565002eec833581210346750032e889c597500000e78020391305816197000000e780e05e2ae613050165ac1b97000000e7802073080c9305016597000000e78020628335012241456394a53a03350121834585002ee2834495008345a500aef98345b500aef58345c500aef18345d5002ef98345e5002ef58345f5002ef183450500aefd83451500aeed83452500aee983453500aee583454500aee1834555002eed834565002ee983358121034a750089c597500000e780002f1305016597000000e780c0542afd1305016597000000e780805e2a8d080c13060002ee8597600000e78040d30345012101c503441121d1aa8335812113852500636eb52a130460036311ad1c4a752205aa75c2050a7662066a682208ca68c208620a939284004e7342032e7462048e76b363d500d18d6e6e220ece66c2062e6762070e65b367a800b3641a01126533e5a20033646400b3e575006e763366ce00d98ec58f418d8215558e8217b3e8a50033e8c7000346811085428347810b6315560a62762206c276c206a274e2048273a20362634203c26ee20e667f220f467e420e267a620a0675b36fa600c58ee660a200466d420da665e205066533e7a30033e66e002a653364af003365ca01b3e6f6018a64b3e49000b3e5a501598e418d8216c58d0216c98e4d8e639857043337c800ba876384d800b3b7d8006395071c3275f265638aa50e3275f265c5a817d5ffff1305c59497d5ffff938645999305b002130601652db1639457083275f2656380a5023275f26531a83275f2656383a5043275f26589a01145f2656ff0af9d1275d26533b6a500631d0616127652673335c700b275f266b385b640898d3305c740b3c5b8003345a8004d8d1304700329e56da01275d2653337b500631907141277d26433359700b275f2679d8d898d33059740b58d318d4d8d1304a00311ed32756386a80032753335150121a01275333505011304800335c10335016597500000e780c0950335816197500000e7800095628597500000e78060945e8597500000e780c093a5b41275d265b3b7a500ede73385d840198db305c84012775266b334e600b276f267b386d740858e198e358db18d4d8d1304900345f10335016597500000e780a08f0335816197500000e780e08e628597500000e780408e5e8597500000e780a08d014411b417c5ffff1305e57f97c5ffff93866504f9bc17c5ffff1305c57e97c5ffff9386c5099305b00213060163e9b417c5ffff1305257d97c5ffff938625084dbc17c5ffff1305057c97c5ffff9386050745b417c5ffff1305e5599305b0026ff02f8b17c5ffff1305e500c9ba17c5ffff130545026ff08f8917c5ffff130585016ff0cf8817c5ffff1305c5006ff00f8817c5ffff130505006ff04f8741456ff0ef8297300000e780a0550000172300006700635f173300006700239c797106f422f026ec4ae84ee43284ae892a89328597200000e780205daa8405c163e38900a2892685ca854e8697600000e78040374a8597300000e78040982685a2700274e2644269a26945618280011106ec22e826e42a8497200000e780e058aa8401c926858145228697600000e78080262685e2604264a26405618280411106e497400000e780c0d90000411106e497400000e780e0d80000397106fc22f82a840a85194697500000e780c0a802650dc14265a26502662af42ef032ec2c08228597500000e78020cee27042742161828017c5ffff1305256797c5ffff938625f29305b002300897400000e780a0d10000397106fc22f82a840a851d4697500000e78040a302650dc14265a26502662af42ef032ec2c08228597500000e780a0c8e27042742161828017c5ffff1305a56197c5ffff9386a5ec9305b002300897400000e78020cc0000397106fc22f82a840a85214697500000e780c09d02650dc14265a26502662af42ef032ec2c08228597500000e78020c3e27042742161828017c5ffff1305255c97c5ffff938625e79305b002300897400000e780a0c60000397106fc22f82a840a85354697500000e780409802650dc14265a26502662af42ef032ec2c08228597500000e780a0bde27042742161828017c5ffff1305a55697c5ffff9386a5e19305b002300897400000e78020c10000397106fcaa852800014697500000e780e092226519cd6265c26522662af82ef432f0081097500000e78080b0e2702161828017c5ffff1305855197c5ffff938685dc9305b002101097400000e78000bc0000397106fc22f82a840a85054697500000e780a08d02650dc14265a26502662af42ef032ec2c08228597500000e78000b3e27042742161828017c5ffff1305054c97c5ffff938605d79305b002300897400000e78080b60000397106fcaa852800094697500000e7804088226519cd6265c26522662af82ef432f0081097500000e780609ee2702161828017c5ffff1305e54697c5ffff9386e5d19305b002101097400000e78060b10000397106fc22f82a840a85154697500000e780008302650dc14265a26502662af42ef032ec2c08228597500000e78060a8e27042742161828017c5ffff1305654197c5ffff938665cc9305b002300897400000e780e0ab0000797106f422f02a840a85194697400000e780807d026519c94265a265026608e80ce410e0a27002744561828017c5ffff1305a53c97c5ffff9386a5c79305b0021306f10197400000e78000a70000011106ec22e826e44ae02e892a84130505041306800b814597600000e780e0f117c5ffff930505c613060004228597600000e78060fd13053900a14522868346e5ff0347d5ff8347f5ff83440500a206d98ec207e204c58f0347150083442500dd8e834735000217a214458fc217830445005d8f1c62d98ee214c58ebd8e14e2fd1521062105c5fd0345090068f4e2604264a26402690561828069ce797106f422f026ec4ae84ee452e03284ae842a89687193050008b389a54063f6c9082330090e130a09065295a6854e8697600000e78060380335090493050508033689042330b904133505f81345150032952334a9044a85d28597000000e78000083304344113051008ce94636fa402930900080335090493050508033689042330b904133505f81345150032952334a9044a85a68597000000e7804004130404f893840408e3e789fc0335090e4a9513050506a685228697600000e780e02f0335090e22952330a90ea2700274e2644269a269026a45618280417186f7a2f3a6efcaebcee7d2e356ff5afb5ef762f366ef6aeb6ee72e892a842801130600082401814597600000e78060d90d0941458345e9ff0346d9ff8346f9ff03470900a205d18dc206620703461900d98e03472900d58d0216834639002217598e03074900c216558ed18d6217d98d8ce07d15a104210955fd280213060004a28597600000e780a0e02c603064833204053267b2772a65aae89776000083b46642033884053e972a97a58db98d9774000083b4a44193d605028215d58d338e9500b346fe004a652ae193d78601a216dd8e2a973303d700b345b30013d70501c215b3e8e500469eb345de0093d6f50386055267d274ea67bee4177500000335653db3ebd50026973e97318d398d9775000083b5a53c135605020215518daa95ad8c8a7636f813d68401a214d18c3386e600330996003345a900935605014215b36cd500338abc0033459a009355f5030605f26672772a769774000083b48438b369b500ba96b296328c32f433c59200358d9774000083b464379357050202155d8daa94258fca752eec935787012217d98fae96b382f60033c5a200935605014215b36dd500ee94a58f13d5f703860792761666ea75aefc177700000337873333eba700b296ae963345e800358d177700000337a7329355050202154d8d2a97398e8e67bef0935586012216d18dbe96b383b60033c5a300135605014215518d2a97b98dae6a13d6f5038605d18d56934e933345a300135605020215498eb29433c53401ce69935685012215c98e338569004ee8b30ed50033c6ce00935706014216336df600b3009d0033c6d0006e6f9356f6030606b36fd6007a99fae033032b01b347130193d407028217c58f3e97b34467010e75aaf493d88401a21433e61401b3086500b298b3c7f80093d40701c21733e39700330be3003346cb002e75aaf81357f6030606b364e600aa92ae9233c69201135706020216598e329eb345be004e7913d78501a2154d8fb30559004af03388e5003346c800935206014216b36256003386c201318fee751355f7030607336ea700ae93ae86aeecde9333c5b301935d050202153365b501b30c4501b3cd7c01926793d58d01a21db3e5bd00be933e873efcb38db30033c5ad00935305014215336a750033059a01a98d93d7f5038605dd8db69eae9eb3c76e0093d607028217dd8e3696b18d93d78501a215dd8db387ee01b38eb700b3c6de0093d70601c216b3e3f6003383c300b345b30013d6f5038605b3ecc500e298fe98b3c5120113d605028215d18d2e953346f501935686012216d18e56e4338658013696b18d93d70501c215b3e8f500b382a80033c5d2009355f50306054d8d4e982698b3450a0193d605028215cd8eb690b3c5900093d78501a215cd8fb3050701b38ff500b3c6df0093d40601c21633e89600c290b3c6f00093d7f6038606d58fca9df29db3c6ad0193d406028216d58c338f6401b346cf0113d78601a216558fe676ee96338ae600b3449a0093d50401c214c58d2e9f3347ef009354f7030607d98c8a66b69eaa9eb3c5be0013d705028215d98d33871500398d935685012215c98e467b33856e01b30ed500b3c5be0013d50501c215b3eba500338deb00b346dd0013d5f6038606b3e0a600466c62963e96334576009355050202154d8d2a9fb345ff0093d68501a215d58d266e7296b309b60033c5a900935605014215558d2a9fb345bf0093d6f5038605b3edd5002676b29fa69fb3c51f0193d605028215cd8e3693b345930093d48501a215cd8c8675fe95b3839500b3c6d30093d70601c216d58f3e93b346930093d4f6038606b3e8960062673a9a669ab3460a0193d406028216c58eb692b3c4920193d58401a214c58d4279b3044901b38fb400b3c6df0093d40601c21633ea9600b3045a00a58d93d6f5038605d58db29eae9e33c5ae00935605020215c98eb382660033c5b200935585012215c98d33855e01b30cb500b3c6dc0013d50601c216b3eea600f69233c5b2009355f50306053363b50033063b010696b18f13d5070282175d8d3388a400b345180093d68501a215d58d62962e96318d935605014215b360d50006983345b8009355f50306054d8dba93ee93b3457a0093d605028215cd8eb387a601b3c5b70113d78501a215b3e4e500b385c301338a9500b346da0013d70601c216b3e3e6009e97bd8c93d6f4038604c58ee275ae9fc69fb3c47f0113d704028214458f3a9fb3441f0193d58401a214c58d827bde9fae9f33c7ef00935407014217458f3a9fb345bf0093d4f503860533ec95008665ae9caa9c33c7ec00935407020217458fba973d8d935485012215c98ce669338599012695298f935807014217336b1701b30cfb0033c79c009357f7030607b36df700ca8a4a96b305d60033c7be009357070202175d8fb307ef00bd8e93d48601a216c58e66762e96338dc6003346ed00135706014216b36ee600338efe00b346de0013d7f603860633efe6000676329a629a33471a00935407020217458fba92b3c5820193d48501a215cd8c8a68b3854801338a95003347ea00935707014217336cf700e292b3c7920093d4f7038607b3e097004267ba9f9a9fb3c77f0093d407028217c58f3e98b344680093d68401a214c58e2279ca9fb69fb3c7ff0093d50701c217dd8db3870501bd8e93d4f6038606c58e329536953346d501935406020216458e33085600b346d80093d48601a216c58e3a953695298e935406014216336396001a983346d8009356f6030606b362d600569d6e9d3346ac01935606020216d18eb69733c6b701135786012216598e3387a801b30ac700b3c6da0093d40601c216b3e39600b38df30033c6cd009356f6030606558e5e9a7a9ab3c5450193d605028215cd8eb3889601b3c5e80193d78501a215cd8fc675d295338ab700b346da0093d40601c21633ef9600fa98b3c7f80093d4f7038607c58fa675ae9f869fb3c66f0193d406028216d58cb38ec401b3c61e0093d58601a216d58db3863f01b38fb600b3c49f0093d60401c214c58eb69eb3c5be0093d4f5038605c58da66b5e953307c500b98e93d406028216c58eb69833c6c800935486012216458e66753a953295a98e93d40601c21633ec9600b30c1c0133c6cc009356f6030606336ed600e26833871a013e9733466700935606020216558e3303d601b346f30093d78601a216dd8e866a5697330dd7003346cd00135706014216598e3293b346d30013d7f6038606b3e0e600ca894a9a2e9ab3467a0013d706028216d98e3698b345b80013d78501a215d98dc66433079a00b38ee500b3c6de0093d70601c216dd8e3698b345b80093d7f5038605b3e3f5006279ca9f969fb3c5ef0193d705028215cd8fbe9db3c55d0013d78501a2154d8f226bb305fb01338fe500b347ff0093d50701c217dd8dae9d33c7ed009357f70306075d8fc2673e953a95298e9357060202165d8e32983347e8009357870122175d8f2695b307e5003d8e135506014216b362a60016983345e8001356f5030605518d2ae8469d729d33c5a601135605020215498eb29d33c5cd01935685012215c98e06756a95330dd5003346cd00135706014216b36fe600338ebf013346de009356f6030606d18ede9e869eb3c5d50113d605028215d18db388950133c61800135786012216598e33873e01b30dc700b3c5bd0093d40501c215b3ee9500f698b3c5c80013d6f50386054d8e569f1e9fb3458f0193d405028215cd8c2693b345730013d58501a2154d8db3052f01b383a500b3c4930093d50401c214c58db3846500258d1357f5030605498f6665aa97b697bd8d13d5050282154d8daa98b3c5d80093d68501a215d58d8a66be96b380b60033c5a000935705014215336af500b30b1a0133c5bb009355f50306053363b50026794a9d329d33c5a201935505020215c98db388b40033c5c800135685012215498e467c33058d01330fc500b345bf0093d70501c215cd8fbe98b3c5c80013d6f5038605b3e2c500667dea9dba9db3c5fd0113d605028215d18d2e983346e800135786012216518f33866d01da89b30ce600b3c5bc0093d40501c215c58d2e983347e8009354f7030607b36f9700c27dee934265aa9333c7d301935407020217d98cb38ac40133c7aa00135587012217598d027e33077e00b30ea700b3c49e0013d60401c214d18c33865401318d9356f5030605558da666b690aa90b3c6f00093d706028216dd8eb38a060133c5aa009357850122155d8db3878001aa97bd8e13d70601c21633e8e600c29a33c5aa009356f5030605b363d5006a9f1a9f33c5e501935505020215c98d2e9633456600935685012215c98e06657a95330dd500b345bd0013d70501c21533e3e500330fc300b345df0013d6f5038605d18d4665aa9c969c33c69401935606020216558eb29bb3c65b0013d78601a216558fb3862c013309d7003346c900935406014216336b9600da9b33c6eb001357f6030606598ece9efe9e33c74e01935407020217d98ca69833c7f801935687012217d98e3387be01330cd700b3449c0013d70401c214458fb3041701a58e13d5f6038606c98e2275aa97ae973d8f135507020217598db30f7501b3c5bf0013d78501a215d98df297338ab7003345aa00135705014215b362e500969f33c5bf008e689355f5030605b369b500469d329d33450d019355050202154d8db30e950033c6ce00ca7d135786012216598eb384ad01338dc4003345ad00135705014215498fba9e33c6ce00926c9357f6030606b36bf60066993699334669009357060202165d8eb29ab3c6da0093d78601a216dd8ee667ca97338ed7003346ce00135506014216518daa9a33c6da009356f60306063369d6008a652e9c1e9c33468b01935606020216d18e369f33467f004e68935786012216d18f33060c01338bc700b346db0013d60601c216558eb306e601b58fae7493d5f7038607dd8dd294ae94258f9357070202175d8f330f5701b3c5e50193d78501a215cd8fb385b401338cb70033478701935407014217336a9700529f33c7e701ca679354f703060733639700ea97ce973d8d135705020215598db303d500b3c6790013d78601a216558fb3869701b30cd70033459501935705014215b369f500ce93334577006e779357f50306055d8d72975e97398e9357060202165d8eb29fb3c7fb014e7e93d48701a217c58f7297338de7003346a601135706014216b36ae600d69f33c6f7012a779357f60306065d8e5a974a97b3c5e20093d705028215cd8fbe9eb345d901ee6693d48501a215cd8cb305d700b382b400b3c7570093d60701c217dd8eb69e33c7d401aa679354f7030607d98ce297aa97bd8e13d706028216d98eb69f3345f501135785012215598dc697330cf500b3c6860113d70601c21633e9e6004ae3ca9f3345f501ea761357f5030605b36be500e696b2963345da00135705020215598d330ad501334646018a7e135786012216598ef696b30dd6003345b501935605014215558d2a9a334646019356f6030606336bd600429d269d33c6a901935606020216558e329fb3c6e401ea6493d58601a216d58db3069d00b38cd50033469601935406014216458e329fb3c5e501ae6493d7f5038605b3e9f500a6929a92b3c55a0093d705028215cd8fbe93b34573008e7493d68501a215cd8eb3859200b38ab600b3c7570193d50701c217dd8db3877500bd8e13d7f6038606d98e629e369e3345c501135705020215598db302e501b3c6560013d78601a216d98e269e338cc60133458501135705014215b363e5009e9233c556009356f5030605336fd5007af6ee98de9833451601135605020215518d3303f50033c66b00ee76135786012216598ec696b30bd60033457501935605014215336ed5007293334566002e769356f5030605558d66965a96b18d93d605028215d58db386f5013347db00ca67935487012217d98c3e96338bc400b3c5650113d60501c215b3efc500fe96b58c93d5f4038604b3ecb400d69ece9eb345d90113d605028215d18d2e9a33c64901935486012216d18c33860e01b38ac400b3c5550113d60501c215d18d2e9a33c64401ca741357f6030606598ee294aa94a58d13d705028215d98dae96358d2a679357850122155d8d2697330de500b3c5a50113d70501c215b3eee50076e3b388de0033451501126c9356f50306053369d500e29be69b33c57301935605020215c98eb383460133c57c002a77935785012215c98f3385eb00338aa700b3c6460113d70601c216558fba93b3c677002e6893d7f6038606b3ebf600429b329bb3466e0193d706028216d58fbe9233465600ea75935686012216558eb306bb00330bd600b3c7670113d50701c2175d8daa92334656006a6e9357f6030606b369f600f29afa9a33c65f01935706020216d18f3e9333466f00ee66935486012216d18c3386da002696b18f93d60701c217dd8e3693b3c7640093d4f7038607c58fea95be952d8f935407020217d98ca69233c75700935787012217d98fe295b38ab700b3c4540193d50401c214b3efb400fe92b3c5570093d7f503ee74860533eff5007af6d294ca94258d935505020215c98d2e9333456900ce67135785012215498f3385f400330ca700b3c5850193d70501c21533eaf5005293b34567000e7793d7f5038605cd8f5a975e97b98e93d506028216d58dae98b3c61b018a7413d58601a216558d2697b304e500a58d93d60501c21533e9d500ca9833451501aa659356f5030605558db295ce9533c6be00935606020216558eb293b3c6790013d78601a216d98ec2953388b60033460601135706014216598eb293b3c676002e7793d5f6038606d58d56973e97398e935606020216558eb298b3c6170193d78601a216d58fb306c701b389d70033463601135706014216b36ee60076e3f69833c617014e779357f6030606336bf60062972a9733c6ef00935706020216d18fbe93334575008e6f135685012215518d3306f701330cc500b3c7870113d70701c2175d8fba93334575004a6e9357f5030605b36af500f294ae9433459a009357050202155d8daa92b3c555002a7a13d68501a215d18dd294b38c950033459501135605014215336dc500ea92b3c555006e6693d6f5038605b3ebd50032987a98b345090193d605028215cd8eb3846600b3459f004a7393d78501a215cd8fb30568003389b700b3c6260193d50601c216d58dae94a58f93d6f7038607dd8e4e963696318f9357070202175d8f33085700b3c60601ea6713d58601a216558d3e96b30dc5003347b701135607014217b369c7004e98334505011356f5032e670605336fc5007af662975a973345ed00135605020215518db302950033465b009357860122165d8e5297330be60033456501135705014215336ae500d292334556001356f5030605518de69fd69fb3c5f50113d605028215d18d3387150133c6ea00ea74935786012216d18f33869f00b38fc700b3c5f50193d40501c215b3e895004697b98f93d5f7038607dd8d4a9e5e9eb3c7ce0193d407028217c58fbe93b3c47b0013d68401a214458e7293b30e6600b3c7d70193d40701c217c58fbe933346760092649356f6030606558eee94aa94a58f93d607028217dd8e3383e600334565000e779357850122155d8d2697b30be500b3c6760193d70601c21633eef60072e3729333456500ce669357f50306053369f500da96ae9633c5d900935705020215c98fbe9333c57500ee75935485012215c98c3385b600338ba400b3c7670193d50701c217dd8dae93b3c674008a7a93d7f6038606b3e9f600d69fb29fb346fa0193d706028216dd8e369833460601ae77935486012216458efe97330cf600b3c6860193d40601c216c58e369833460601ce741355f6030606336aa600a69efa9e33c5d801135605020215518daa9233465f002a67935486012216458eba9e330fd6013345e5019357050142155d8daa92334656009357f60306065d8e5e973297b98d93d705028215dd8d2e9833460601ca67935486012216d18c3306f700b38cc400b3c5950113d70501c215b3efe5007e98b3c5040113d7f503ea678605b3eee50076f6da97ca97bd8e93d506028216cd8eb3885600b345190113d78501a2154d8fb3855701330bb700b3c6660193d70601c216b3eaf600d69833471701aa779354f7030607458fe297ce973d8d935405020215458d2a93b3c46900ca7693d58401a214c58dbe96b38bd500334575019356050142153369d5004a9333c56500ea759356f5030605c98efa95d2953345be00935405020215c98ca69333457a008e67135685012215498e3385f500330ca600b3c4840193d50401c214c58db38775003d8eae629354f6030606458e969cba9cb3c5950193d405028215c58db3836500334777004e63935487012217458fb3846c00330d9700b3c5a50113d50501c21533efa500fa9333457700ee6c9355f5030605b369b500669b369b33c56f019355050202154d8daa97bd8e8e7513d78601a216d98eda95338bb60033456501135705014215498f330ef70033c5c601ae769357f5030605336af500de96b29633c5da009357050202155d8d2a9833460601ce7f935786012216d18f3386f601b38bc70033457501935605014215558d2a98b3c50701ee7793d6f5038605b3ead5003e9c769cb345890193d605028215d58dae98b3c41e01926613d68401a214458eb304dc0033099600b3c5250193d40501c215c58dae98334616019354f6030606458eea97b2973d8f935407020217458f3a9833460601935486012216458ee697330cf60033478701935407014217b36e97007698334606011357f6030606aa74598e7ae332f6da94ce94258d135605020215518d3306150133c7c900935787012217d98f33875400b389e70033453501935405014215b36895004696b2ea3d8e1355f6030606b367a6005e93529333c565009355050202154d8daa93b3457a0013d68501a215d18d3306d3003383c50033456500935605014215b362d500969333c575009355f5030605b366b500ca9fd69f3345ff01935505020215c98d2e9e33c5ca01ea74135685012215498e33859f00330fa600b3c5e50193d40501c215cd8c269eb345c6014a6613d5f5038605c98d62963e96b18c13d504028214458daa93b3c77700ae7413d78701a2175d8f26963a9632e6318d135605014215518d2ae31e95aaee398d1356f5032a670605518d2afa4e97369733c5ee00135605020215518d2a9e33c6c601ea669357860122165d8eba96b29636ea358d935605014215558daaf67295aaf2318d1356f5038e760605518d2afe9a96ae9633c5d800135605020215518d2a98b3c505010e6613d78501a215d98d36962e9632ee318d135605014215518daafa4295aae62d8d9355f50306054d8daae23275ca75aa95fa9533c6b200d666135706020216598eb296358d0a779357850122155d8dba95aa952ef2b18d13d60501c215d18daefeb695aeea2d8d9355f5030605c98da8022ef6a1451060833605fc1861358e398e10e0fd1521052104f5f5be701e74fe645e69be691e6afa7a5a7bba7b1a7cfa6c5a6dba6d7d618280197186fca2f8a6f4caf0ceecd2e8d6e4dae05efc62f866f46af06eec906103bc8500329c636fcc34aa8988699376f50093b616003337a000f98e6380063a814a89466368d5008d462a87850a0581e3ede6fe83cb85013285d68597000000e780a03b6365ac322a8d1305000463f5aa323305ac4133555501814c89456368b5008d452a86850c0581e3edc5fe938d2c0063ea9d316145b3b5ad02639a0530b384ad02ea9463eaa43113893c006a847d19268a630d0902630c0d24233044015285639b0b00130600105285814597400000e78060200860610408e1c10408e5e3f844fd17a5ffff13052506a5ac4ee0638b0d2e014b13098d0093891c005a85ee8597000000e780a03563030d201d05935435002330490163990b0052858145268697400000e780201bd29463e24425638669016109050b268ad1b7094963e72d0593098d02330a904105442285ee8597000000e780c0301d05135b350023b0990063990b00268581455a8697400000e780801633856401636195200504b3058a00e109aa84e39325fd11a02685d68597000000e7806028636fac2463860d262a8b938bfdff2a84638b0b161385edff9305f00363eda520854c5a846ae86ee463080d14aa843395ac00331d55013309a401636589186145b38da402c265ae9d3385ab022e9593098500130a0501636f2c0d03b50d000c612300b40013d68503a303c40013d605032303c40013d68502a302c40013d605022302c40013d68501a301c40013d605012301c400a181a300b40093558503a307b400935505032307b40093558502a306b400935505022306b40093558501a305b400935505012305b40093558500a304b4002304a4000c6180e500e15a85d6852686a28697000000e780c022058915ed5a85d6855e86a28697000000e780802183b5090013563500b295838605001d893395ac00c98e2380d50083350a00b29503860500518d2380a5004a846a99e37489f249a82685a26597000000e780c0185a85d6852686a28697000000e780801c83b58d0013563500b295038605001d893395ac00518d2380a50081cc1385f4ffa68b426de31c0dea97200000e78020b00000426da26d63638c0a33058c40826523b0650123b4850188e923bca50123b0b50323b45503e6704674a6740679e669466aa66a066be27b427ca27c027de26d0961828017a5ffff1305a5def14597200000e780e08e000017a5ffff130565ddf5b717a5ffff1305c5dccdb717a5ffff130525dce1bf17a5ffff130585d5ada817a5ffff1305e5d793054002c9b717a5ffff130505da5dbf17a5ffff130565d0a1a817a5ffff1305c5d84db717a5ffff130525d291a017a5ffff130585cb9305300271b717a5ffff1305a5da29a85285d68597000000e780c002637bac0017a5ffff130585dd97000000e7804005000017a5ffff1305e5cd9305100289bf01cd1306000463f0c5027d153355b50005053315b500828017a5ffff130585cb9305100239a017a5ffff1305a5cd9305400297200000e780c080000097200000e780e09c000063efa5006382a5021345f5ffaa951305000463f2a50205453315b500828017a5ffff1305c5c629a017a5ffff130525c69305100239a017a5ffff130545bf9305300297100000e780607b000063e0a6041307f003636cc7001307000463fde500898e33d5c6003355b500828017a5ffff1305e5c429a017a5ffff130545c49305400297100000e7806077000017a5ffff130565cfb545f5b790659461137806fc3698636bd80c98699355660063e3e500ba8594e2094694e6b68763ebc508fd1593d8860393d2060313d3860293d3060213de860193de060113df8600b68736863e879387070463efe7062380c70013578603a383e700135706032383e70013578602a382e700135706022382e70013578601a381e700135706012381e7002182a380c7002384d700a387170123875700a386670023867700a385c7012385d701a384e70190621ce6fd159ce23e86c9f99385070463e7f50214e1233405010ce914ed828017a5ffff130565b8f14597100000e780a068000017a5ffff130525b7f5b717a5ffff130585b6cdb7717106f522f126ed4ae94ee552e1d6fcdaf8def4e2f0e6eceae82a841305000497550000138ae5436371850417550000930425438860631e05348864fd558ce063130512c870cc6cd068d464aae4aee032fc36f80a850c1897000000e780209c054588e413850401c5a803350a04631b053203358a04fd552330ba041ded03350a0883358a0703360a07aae02efc32f80a850c1897000000e78080e705452334aa040265a2654266e2662338aa04233cba042330ca062334da0603398a0663000902033509000c6110650ce20c6510610ce6130b0a04630825032a8991a403390a0603358a056373a902130509046368252983350a042330aa0685052330ba046315092209a823340a0619ac03350a0405052330aa0403350a00631e052803358a00fd552330ba001ded03350a0a83358a0903360a0983368a08aae4aee032fc36f80a850c1897000000e780408d05452334aa0013050a018a851306000397400000e780c0c583398a031305f003636335210545814c3315350163788500850c63840c1c0605e36c85fe83350a0363e3bc00e68503358a020146e146b386dc02aa96138406fdb385bc406389c516630d051c147803b9060061047d16e307d9fe033509008335890088e1033589008335090088e5047017550000130b852803350b0183358b03934af6ffe69a5686ca8697000000e78000cd93553500a695038605001d89854b3395ab00518d2380a50063f85c11130c000417550000130b6524138afaff63778a1333954b01b3143501ca9463e72413033d840203350b0183358b035686ca8697000000e780a0c793553500ea95038605001d893395ab00518d2380a500833a840003350b0183358b035286ca8697000000e780c0c493553500d695038605001d893395ab00518d2380a50008600c612380b40013d68503a383c40013d605032383c40013d68502a382c40013d605022382c40013d68501a381c40013d605012381c400a181a380b40093558503a387b400935505032387b40093558502a386b400935505022386b40093558501a385b400935505012385b40093558500a384b4002384a4000c6184e504e12114d28ae3e54cf119a00149528b03350b0005052330ab004a85aa700a74ea644a69aa690a6ae67a467ba67b067ce66c466d4d61828017a5ffff1305658121a81795ffff1305c5749305300231a01795ffff1305e57ff14597100000e780203000001795ffff1305a572f9bf1795ffff1305057ecdb797100000e780204a000017a5ffff1305d5b49795ffff9386c56d15a017a5ffff1305b5b39795ffff9386a56c09a817a5ffff130595b29795ffff9386856bc1450a8697100000e78020450000317106fd22f926f54af14eed52e956e55ae1defce2f8e6f4eaf0eeec97550000938ce50683b50c04639d05382a8903b58c04fd5523b0bc041de9175500001304050548602c7c3078aae4aee032fc28002c1897000000e78060ae054528e42265c2656266827628e82cec30f034f403b50c0583b58c053335a9001345f5ffb335b9006d8d51c517550000130545002c75638e052090612300c90093568603a303d900935606032303d90093568602a302d900935606022302d90093568601a301d900935606012301d9002182a300c90013d68503a307c90013d605032307c90013d68502a306c90013d605022306c90013d68501a305c90013d605012305c90013d68500a304c9002304b900906165a203b50c0483b50c00050523b0ac04639b052a03b58c00fd5523b0bc0015ed175500001304c5f548704c6c50685464aae8aee4b2e036fc28002c1897f0ffffe780c04f054508e4130504012c001306000397400000e780608883ba0c03638f0a2283b98c02138afaff13848902854463809a04638b0922033b040003b50c0183b58c032686ca8697000000e780609593553500da9583c505001d8933d5a50005898504610469d5f91463e6440139a263030a108144930a0004268b63e49a00130b000483bb8c0303bc0c0161453385a4024e9513048502054d03b50c0183b58c032686ca8697000000e780808f638e091a833504fe13563500b2950386050093767500b316dd0093c6f6ff758e2380c500937515003306b040833604fe13661600329513563500369603460600937675003356d600058a51e2630b9b1263fe5b1333159500331575016295636e85131061146590e21065146190e691c12a89833d040003b50c0183b58c0385042686ca8697000000e780c08693553500ee95038605001d893315ad001345f5ff718d2380a5006104e3129af4d28405a023302901930585064a862334260123b02501930c050451a8638a090e814461453385a4024e9508610c612300b90013d68503a303c90013d605032303c90013d68502a302c90013d605022302c90013d68501a301c90013d605012301c900a181a300b90093558503a307b900935505032307b90093558502a306b900935505022306b90093558501a305b900935505012305b90093558500a304b9002304a9000c6123b425012330250103b50c00050523b0ac00ea704a74aa740a79ea694a6aaa6a0a6be67b467ca67c067de66d296182801795ffff1305c53429a01795ffff130525349305300231a01795ffff1305453ff14597100000e78080ef00001795ffff1305053893051002edb797100000e780e00900001795ffff130595749795ffff9386852d09a81795ffff130575739795ffff9386652cc145300097100000e780000600005d7186e4a2e026fc4af84ef452f056ec83ba050263800a0a2e8a2a898065b35954034e8597000000e780200b83340a002ae02ee402e863e335078145636e54031396350032950d466370560983c6140003c70400a206d98e03c7240083c7340033045441d6944207e2075d8fd98e14e185052105e37a54fd2ee8226502662338b9002334a9002330c900a6600664e2744279a279027ae26a616182800a8581454e8697000000e7806008c2650265e37954f9d9b71795ffff13054539e54597100000e78080de00001145d68597100000e780e0570000011106ec22e826e42a841dc51355c40305ed93351500931434008e0599c4268597200000e780800eaa8581e9268597200000e780a00f0000a1452e85a285e2604264a2640561828097d0ffffe780401b0000411106e497000000e78000037d567e1605066315c500a2604101828011e597d0ffffe780c01800002e8597200000e780c00a00005d7186e4a2e026fcae86b29563f4d5000145a1a82a8408659314150063e39500ae84914563e39500914493d5c40393b51500139634008e0501c914600e0536f0a14636f42af811a002f42800141097100000e780606aa265426599c1e26531a008e004e47d557e150505a6600664e27461618280411106e4054697000000e78060f87d567e1605066315c500a2604101828011e597d0ffffe780200e00002e8597200000e78020000000797106f422f026ec4ae84ee452e06365d7046366e604aa89b304d7403389d5002685814597100000e780806b2a842e8aca85268697300000e780a03b23b0890023b4490123b89900a2700274e2644269a269026a456182803685ba8519a03a85b28597100000e780203e0000797106f422f026ec4ae84ee452e06363d604aa89b304d6403389d5002685814597100000e78000652a842e8aca85268697300000e780203523b0890023b4490123b89900a2700274e2644269a269026a456182803685b28597100000e7800038000063e8c60063e9d500b385c640329582803285b68511a0368597100000e780e0350000011106ec22e826e42a8410690865ae846319a6002285b28597000000e78020ec10680860931536002e9504e1050610e8e2604264a26405618280397106fc22f826f44af04eec52e856e4114a32892a84637d46032d45ad4a814597100000e7802059aa84ae891795ffff9305e5132d46268597300000e780c028054508c0233444012338240104ecb1a803c5150003c6050083c6250083c535002205518dc206e205d58db3e4a500b9c09104638424052d45ad4a814597100000e78060532a8aae891795ffff9305250e2d46528597300000e78000232320040004e423382401233c4401233034032334540331a0114a631d4901154508c0e2704274a2740279e269426aa26a216182802d45ad4a814597100000e780c04daa84ae891795ffff930585082d46268597300000e780601d23200400a9b71061833805011c65210605483e8763ee17019307f7ff10e11ce5637d1801833686ff0c622106e3f3d5fe333517011345150082800545854597100000e780601e0000411106e410610e069796ffff938626d2369610620286907588711c6e9795ffff9385950d3d4635a8907588711c6e9795ffff9385c50b2d462da021052ae01795ffff9307c5071795ffff130745083d463da0907588711c6e9795ffff9385a5042146a2604101828721052ae01795ffff9307c5001795ffff1307e5001d468a862e85be8597100000e780000ca2604101828082808365050005466345b60099c9054609a809466389c5000d466394c500210521a0610511a041050c6591c5086117230000670083cb8280397106fc22f83287ae862a8402f002ec02e802e4130500022af405659b0815822c108d472800894201460148730000006309550285456308b502914515e522751306000289456361a602130514002c001306000297300000e78080062300040009a8854511a081450ce408e805452300a400e270427421618280397106fc22f83287ae862a8402f002ec02e802e4130500022af405659b0815822c109547280089420146014873000000630b55028545630cb502914515e922751306000289456365a602130524002c001306000297300000e780e0fe01458545a300b40009a80145a300040029a081450ce408e805452300a400e270427421618280130101ba233c1144233881442334914423302145233c3143233841432334514323306143233c7141b289ae8b2a8408081306004093040040814597300000e78080eb2338914005659b08c58293050141080889440146de864e8781470148730000006301950885456300b508914535ed03390141130500406372250b8545054b4a8597100000e780c0222a8aae8a0c081306004097300000e780c0f2930209c013050a402338514085659b88c58293050141130600408944de864e87814701487300000063019508630e6507114b25ed03350141094b63e8a2062330440123345401b1a8854511a081450ce408e8233004008330814503340145833481440339014483398143033a0143833a8142033b0142833b81411301014682804a85814597100000e780e018aa84ae890c084a8697300000e78000e904e0233434012338240145bf014b2334640108e823300400e3810afa528597200000e780c0a551bf9308d0057d558145014681460147814701487300000001a0086101a08280797106f42e8813564500130f7002130710279796ffff938e26e16363e608130f700213076102174600008338064939661b03068f05669b03b6479302c0f937e6f5051b0ef60faa86333515032d813b066502b307d600139607034992330676029355160141821376e67fbb855502be95769683471600c615c19103460600a30ff7fef69583c7150083c50500711f230fc7fea300f7002300b7007117e365defa130630066370a60493150503c99105661b06b647b385c502c5811306c0f93b86c502329546154191791f7695034615000345050093061100fa96a380c6002380a6002e85a945637cb5009305ffff130611002e961b0505032300a60005a006059305efff7695034615000345050093061100ae96a380c6002380a60093061100ae96130770020d8f1795ffff9305e50b4285014697000000e780e000a27045618280597186f4a2f0a6eccae8cee4d2e056fc5af85ef462f066ec6ae86ee4aa8403654503ba893689328aae8b937c1500b70a110063840c00930ab00293754500ce9c89e5814b8c6085e5a1a08145630e0a005286de86038706008506132707fc134717007d16ba957df6ae9c8c6095c103bd840063ffac01218925ed83c58403054633059d41634cb60af9e1aa8c2e85c9a0807084742285a6855686de86528797000000e7806014054b0dc15a85a6700674e6644669a669066ae27a427ba27b027ce26c426da26d656182809c6c2285ca854e86a6700674e6644669a669066ae27a427ba27b027ce26c426da26d6561828780581305000383c584032ee003bc040283bd840288d8054b238c64036285ee855686de86528797000000e780e00c51f5228a33049d4105047d1451c803b60d02930500036285029665d985bf09466398c50093051500058193dc150011a0814c03bc040203bd84028458130415007d1409c803360d026285a68502966dd9054b2dbf37051100054be389a4f26285ea855686de86528797000000e780e00511fd83368d016285ca854e86829619f5b30990417d5a7d59338529016309450303360d026285a6850296050975d50da083b68d016285ca854e868296e31005ee014b23a844030265238ca402c1bd6689333b9901e1b5797106f422f026ec4ae84ee49b070600370811003a89b6842e84aa896389070114704e85b2858296aa85054591ed81cc1c6c4e85a6854a86a2700274e2644269a269456182870145a2700274e2644269a269456182805d7186e4a2e026fc4af84ef452f056ec5ae85ee483320500146933e7d2003289ae896304072a638706101c6d8146338e29018507370311009308f00d1308000f4e8601a893051600918eae962e866303640efd17adc7630fc60d8305060013f4f50fe3d105fe834516009374f40113f7f50363fa8802834526001a0793f5f503b363b7006367040383453600f614ad909a0393f5f50333e4b300458c630c64089305460055b79305260013946400598c61bf93053600b20433e4930071b7630bc6078305060063d3050493f5f50f1307000e63ede5021307000f63e9e50203471600834726001377f70393f7f70303463600f615ad9132079a075d8f1376f603598ed18d370611006386c50285c263fd2601b385d90083850500130600fc63d7c500814591e539a0e39d26ffce8599c13689ae89638b021803388500930500026372b902814e63060916ca85ce86038606008506132606fc13461600fd15b29efdf581aa13877900619b3386e940b308c90093f678008145630d3701ce87038407008507132404fc934414000506a6957df6014691ce93f788ffba9783840700850793a404fc93c41400fd162696fdf693d638009747000083b7e7f89744000083b2e4f8b714001092048504939804018508b30eb6001da013173e001a97b386c34113763e00b3f45500a181b3f55500a695b3851503c191ae9e2deaddcab6833a839305000c368e63e4b600130e000c9375ce0f139435001a94dddd81451a8745df146393c4f6ff9d8099821067c58efd8eb6959346f6ff9d82046b1982558e7d8e93c6f4ff9d829980c58e046ffd8e3696b29513c6f4ff1d829980458e7d8e13070702b295e31d87fabdb7630803029305000c63e4b3009303000c814593f633008e06106021041347f6ff1d831982598e7d8ee116b295f5f611a0814533f65500a181b3f55500b295b3851503c191ae9e63fc0e01834685030546b305d8416345d60285ce814a25a80c7508719c6dce854a86a6600664e2744279a279027ae26a426ba26b6161828709466398c600138615008581935a160019a0ae8a8145033b0502833b85020459138415007d1409c803b60b025a85a68502966dd9054a81a037051100054a638ca40283b68b015a85ce854a86829605e533095041fd597d5433058900630a350103b60b025a85a6850296050475d511a05684333a54015285a6600664e2744279a279027ae26a426ba26b61618280411106e497000000e780801c0000197186fca2f8a6f4caf0ceecd2e8d6e4dae0b2891306000232f80d46230cc10203b4090202e002e82af02ef461c003b589026307051083b409009305f5ff8e058d8113891500a10493058003330ab5026104854a17050000130b458a906001caa276027583b584ff946e829665ed08482ad803058401230ca1024c4803b509012eda033684ff0c6001ce631756019205aa95906563046601014621a08c618c61054632e02ee4033684fe833504ff01ce631756019205aa95906563046601014621a08c618c61054632e82eec0c6492052e95106508618a85029649e5c104130a8afc13048403e31b0af6b1a003ba890163080a0483b4090103b409001305faff12051181130915002104a104120a106001caa2760275833584ff946e829639e1906003b584ff8a8502960ded4104411ac104e31e0afc03b589006368a9002da0014903b589006371a90203b5090012092a99a27602758335090003368900946e829619c1054511a00145e6704674a6740679e669466aa66a066b09618280907588711c6e9785ffff9385b5532d468287907588711c6e9785ffff9385455339468287411106e497000000e78080010000411106e497000000e780a0000000411106e497c0ffffe780401c0000757106e5014730012948bd4821a89306f6ff13d547009a92a30f56fe0507368663fcf800aa879372f50013030003e3e002ff13037005e1bf13050008198d130610086370c5021785ffff9307e55009462e85be8597000000e7800082aa60496182809305000897000000e78040560000757106e522e1a6fccaf8cef4d2f0d6ecdae8dee4e2e066fc6af86ef432892e8a014c814c81499745000003bba5b69745000083bba5b69745000083b4a5b600690c612ef008652aec13058a002ae01785ffff130525482ae8294d22e40da03305b6000345f5ff5915133515002300a4006265146d02758296ee8c6311051213f5f90f631b051063758901e9a8636c890d33058941b3058a014146637fc50063022c0d81463386d50003460600630da6098506e319d5fe75a013867500937686ff3386b640ad8e93b6160013371600d98ea1c20146930605ff02676297b387c5009c6313c4f7ffa58fda9733747401e18f8defb307c7009c6313c4f7ffa58fda9733747401e18f95e34106e3f9c6fc31a83387d500034707006307a7038506e319d6fe930605ffe3f9c6fa6304c5062264b386c50083c606006386a6010506e319c5fe05a0b286e296138c1600e3f026f5d29603c50600e31ba5f38149e28de28a39a04a8c8549e68dca8a63872c030345040001c96265146d11460275c265829611ed33869a41b3059a01e39a9aed0145f1bd4a8c2264f9b7014511a00545aa600a64e6744679a679067ae66a466ba66b066ce27c427da27d49618280411106e41b8605009306000802c26376d6002302b100054671a01bd6b50019ee13d665001366060c2302c10093f5f50393850508a302b1000946ada01bd6050115e613d6c5001366060e2302c10013964503699213060608a302c10093f5f503938505082303b1000d462da81396b50275921306060f2302c1001396e502699213060608a302c100139645036992130606082303c10093f5f50393850508a303b10011464c0097000000e780e0d9a26041018280397106fc907594712ae032f836f4886d906994658c612af032ec36e82ee41785ffff930525320a85300097000000e780a0b2e27021618280086117030000670063d5411106e408611b8605009306000802c26376d6002302b100054671a01bd6b50019ee13d665001366060c2302c10093f5f50393850508a302b1000946ada01bd6050115e613d6c5001366060e2302c10013964503699213060608a302c10093f5f503938505082303b1000d462da81396b50275921306060f2302c1001396e502699213060608a302c100139645036992130606082303c10093f5f50393850508a303b10011464c0097000000e78060caa26041018280397106fc90759471986d32f836f43af0906994658c61086132ec36e82ee42ae01785ffff930585220a85300097000000e78000a3e27021618280357106ed22e926e54ae1cefcd2f8d6f42a840345050109c5833a04008544d5a0b2892e89033a840003654a03833a04009375450091e93336500163880a021785ffff9305e50f35a063960a0483358a0203350a02946d9785ffff9385850e094682961dc5814a854469a81785ffff9305650d83368a0203350a02946e05068296854441e103b689014a85d28502968da803254a038544a303910283350a0203368a022ee432e8930571022eec83250a0303068a0383360a0003378a0083370a0103388a01aaceaecc2300c10636f43af83efcc2e02800aae403b689011785ffff13052502aae82c104a85029619e9c6652665946d9785ffff9385650409468296aa8423089400850a233054012285ea604a64aa640a69e679467aa67a0d618280397106fc22f826f44af02a841c7508719c6f3a89b684829722e8230ca10002e4a30c01002800a6854a8697000000e78060eb22658345810139c50544b9e5834591017d1513351500c264b335b0006d8d05c103c54403118901ed8c748870946d9785ffff938515fc05460544829611ed8c748870946d9785ffff9385a5f4054682962a8419a03334b0002285e2704274a274027921618280411106e497000000e78040a200001785ffff9306850709462e85b68517f3ffff6700834c397106fc22f826f42e848c752ae40870946d9785ffff938585074546829622ec2300a10202e8a30001021785ffff1306050408082c0097000000e780e0de42658345010239c50544b9e5834511027d1513351500e264b335b0006d8d05c103c54403118901ed8c748870946d9785ffff938595ef05460544829611ed8c748870946d9785ffff938525e8054682962a8419a03334b0002285e2704274a27421618280757106e5014730012948bd4821a89306f6ff13d547009a92a30f56fe0507368663fcf800aa879372f50013030003e3e002ff13037003e1bf13050008198d130610086370c5021785ffff9307e5e709462e85be8597f0ffffe7800019aa60496182809305000897000000e78040ed0000797106f422f026ec4ae84ee42a8404690865ae893309b640058d6363250308602695ce854a8697200000e780e0e4ca9404e8a2700274e2644269a269456182802285a6854a8697000000e780c0000468f9b75d7186e4a2e026fc2e966368b6042a8408659314150063639600b284a14563e39500a14493c5f4fffd9119c5106032f0054632f42af811a002f428001410268697000000e780e003a265426581cdfd55fe158505630ab50009ed97c0ffffe78060aa000008e004e4a6600664e27461618280626597100000e780809b0000011106ec22e826e44ae03289aa8499cd2e84886605c18c6a91cd88624a8697100000e780009805e180e419a023b40400854521a8630409024a85a28597100000e780209575d1814588e423b824018ce0e2604264a264026905618280228565f5e1b703e6450308619376060189ea1376060219ea086117f3ffff6700c3ee086117f3ffff6700037b086117030000670063e3411106e422e02a8411c96347040289c9228597100000e780209009a8054501a88545228597100000e780808d19c9a285a26002644101828097c0ffffe780809b0000228597100000e780808d0000797106f422f026ec4ae84ee42a8904690865058d2e84636fb50283390900894533859900636cb4007d148145228697200000e78080bca2943385990023000500850423389900a2700274e2644269a269456182804a85a685228697000000e780e0008334090155bf5d7186e4a2e026fc2e966368b6042a8408659314150063639600b284a14563e39500a14493c5f4fffd9119c5106032f0054632f42af811a002f428001410268697000000e780e003a265426581cdfd55fe158505630ab50009ed97c0ffffe780008e000008e004e4a6600664e27461618280626597000000e780207f0000011106ec22e826e43284aa8499cd88660dc18c6a99cd8862228697000000e780e07b19ed85458ce431a823b40400854511a88545228597000000e78020797dd1814588e480e88ce0e2604264a26405618280411106e422e02a8408617d1508e005e90c70086c8c6182950870086511c5086c97000000e780e075087811c5087497000000e780007508647d1508e409c5a2600264410182802285a2600264410117030000670003735d7186e4a2e026fc4af84ef452f056ec83ba0501368a3289aa8963e3da00d28a806108687de1286c7d5610e8637c55010870106c98651c6d4e85b2854a86d286829761a08465306463edc400b386540163ee96082c683307b600636ec7086376d70208700c6c1074147c1c6d0a85268782970345010069e9a26563e8550f286c2ce824e426866367b50eb3b6c400918c33359500558d49e5338554016363950463e7a5080c7c63eca508b3059540639745090c74a6954a85528697200000e780c0a723b45901238009000868050508e8a6600664e2744279a279027ae26a616182801785ffff130585c311a81785ffff1305e5c229a01785ffff130545c2f14597f0ffffe780802e00001785ffff130515b59785ffff938605b6c1450a8689a01785ffff130505c69305f002d1bf1785ffff130515c893052003d9b7528597000000e780e0a400001785ffff130525d99785ffff9386a5ba9305b0021306710197f0ffffe780804300001785ffff1305c5bc71b71785ffff1305e5bd9305e00241b7034505000e051786ffff1306a6e12a969786ffff938606e6369598751062146188711c6fb6858287411110650c69b29563edc50008611069fd568582637dd60028616369b502410182801785ffff13056589a14535a01785ffff1305a5ab9785ffff9386a5ace145300097f0ffffe780c03a00001785ffff1305b5be9305600297f0ffffe780601e0000797106f422f0aa8502c2280050009146114497000000e78020de0345810011e942656319850203654100a2700274456182801785ffff1305c5c99785ffff938645ab9305b0021306f10197f0ffffe780203400001785ffff130575bab54597f0ffffe780e0170000797106f422f09c6185079ce19dc7b2962ee463e6c6022a8436e83aec280097000000e78080f16265c265226608e80ce410e0a270027445618280000000001785ffff130585a19305b00297f0ffffe780a0120000197186fca2f8a6f4caf0ceecd2e8d6e4dae05efc03bb050003370b00846594692a89130517002330ab006dcd5ae409072330eb0065cbb28a36f85af02e8597000000e78060f09385440063ef950caa892ef4081097000000e78000ef8d4563faa50c09811304f5ff63fe8a02938b1a0013952b0026956364950c2af4081097000000e78060ec2a8a63998b0233854401636c950a2ae863f649051785ffff13058596f1a015452304a900233009005a8597000000e78020c3b1a08a0a33859a002105636895082af4081097000000e780a0e7b385440163e39508aa892ee863644509338549412aec280097000000e78080df6265c26522662338a9002334b9002330c9005a8597000000e780c0bde6704674a6740679e669466aa66a066be27b09618280000000001785ffff1305a58d3da81785ffff1305a5a1b9451da81785ffff1305458c25a01785ffff1305a58b39a81785ffff1305058b11a81785ffff1305658a29a01785ffff1305c5899305b00297f0ffffe780e0fa0000397106fc22f826f42a8402e408083000a146a144a28597000000e78060ba0345010105e16265631f9502a264086097000000e78080b32685e2704274a274216182801785ffff130545a59785ffff9386c5869305b0021306710297f0ffffe780a00f00001785ffff1305a597b94597f0ffffe78060f30000397106fc22f826f42a84a307010008081306f10085468544a28597000000e780a0b2034501010de16265631095048304f100086097000000e780a0ab2685e2704274a274216182801785ffff1305659d9775ffff9386e57e9305b0021306710297f0ffffe780c00700001785ffff1305a590b54597f0ffffe78080eb00005d7186e4a2e026fc4af8ae842a898c69054632e002e402e889c90a8597000000e780c0910266426411a001442808a685a28697000000e78040a9034581011de5027563168504c2652266826688602338b9002334c9002330d900a6600664e27442796161170300006700c3a01785ffff130545939775ffff9386c5749305b0021306f10297f0ffffe780a0fd00001785ffff13055587c94597f0ffffe78060e10000011106ec22e826e49c692a84637df700b384e74063e3d400b684b306970063ede60263f7d7001545a300a400054531a8998e639dd4028c61ba953285268697100000e780c051014504e42300a400e2604264a264056182801775ffff1305656ef14597f0ffffe780a0da00002685b68597f0ffffe780005400005d7186e4a2e026fc4af84ef452f02e8483b905012a896145a14597000000e780000b59c1aa84086888e8086488e4086088e0054a52e402e802ec1314ba002800a28597f0ffffe780a07d13050006a14597000000e780a00731c923304501233445012338050004ed9775ffff938545790cf1a2650cf5c2650cf9e2650cfd23303505233405042338050420ed23340900233839012330a900a6600664e2744279a279027a61618280614519a01305000697000000e780a00300000c6591c508611703000067002301828017b3ffff6700630617b3ffff6700630617b3ffff6700630617b3ffff6700c30a97b0ffffe780200e00005d7186e4a2e026fc4af8ae84806590612a892800a28597e0ffffe78040390345810019c5426529e109452300a90029a805040dc09305910080e4130610024a8597100000e780c03aa6600664e2744279616182801775ffff1305c571f14597f0ffffe78000c4000097f0ffffe78020e00000357106ed22e926e54ae1cefcd2f8d6f4daf02e89aa8a2800d68597000000e78040f7034581008944630b951675cd0345210283451102034631028346410222054d8d4206e206558e518d83456102034651028346710203478102a205d18dc2066207d98ed58d82154d8daae40345a101834591010346b1018346c10122054d8d4206e206558e518d8345e1010346d1018346f10103470102a205d18dc2066207d98ed58d82154d8daae00345210183451101034631018346410122054d8d4206e206558e518d83456101034651018346710103478101a205d18dc2066207d98ed58d82154d8d2afc0345a100834591000346b1008346c10022054d8d4206e206558e518d8345e1000346d1008346f10003470101a205d18dc2066207d98ed58d82154d8d2af829a082e482e002fc02f803b58a010c6903b40a0113060002639bc5040c6108181306000297100000e78080650125854421e103b50a0210610818a28597e0ffffe7808025c279638f09120665627bc145637fb50263070b004e8597000000e780c0de8144130550032300a90011a08544050475c823b88a002685ea604a64aa640a69e679467aa67a067b0d6182804145814597f0ffffe780004b2a892e8a4146ce8597100000e780201b0345190083450900034629008346390022054d8d4206e206558e518d83455900034649008346690003477900a205d18dc2066207d98ed58d8215c98d03459900034689008346a9000347b9002205518dc2066207d98e0346d90033e7a6000345c9008346e90022068347f900498ec20603b58a02e207dd8e558e14651c610216598e3696be9533b7f5003a966304d6003337d60015ef0ce110e563070a004a8597000000e780c0cf63070b004e8597000000e780e0ce03b40a0131b71775ffff13052547f14597f0ffffe780609900001775ffff1305e545f5b71775ffff130545479775ffff9386c54b9305b002900897f0ffffe780c0b100000e059775ffff9385a5c72e950c6105458285094582800d4582801145828097f0ffffe78000b10000357106ed22e926e54ae1cefcd2f8d6f4daf02e8a2a8908100546814597e0ffffe780a002034501020dc12275c27597000000e780a0faea604a64aa640a69e679467aa67a067b0d61828003156102831541020356210283461102231ea104c205d18da274627503560104c27aaeccaae42318c104f5c603150105a6652314a1002ee013050002130b0002814597f0ffffe780a02e2a84ae89ac08194697100000e780a04313d58403a306a40013d504032306a40013d58402a305a40013d504022305a40013d58401a304a40013d504012304a40013d58400a303a4002303940013d58a03a30aa40013d50a03230aa40013d58a02a309a40013d50a022309a40013d58a01a308a40013d50a012308a40013d58a00a307a40023075401130564018a85294697100000e78040f68144631c6a01130600022285ca8597100000e78060379334150063870900228597000000e780e0b213057004e38f04ec0145e1bd3945d1bd130101c0233c113e2338813e2334913e2330213f233c313d2338413d2334513d2330613d233c713b93070002631df6503a8ab6892a8903c5950103c6850183c6a50103c7b5012205518dc2066207d98e558d03c6d50183c6c50103c7e50183c7f5012206558e4207e2075d8f598e0216518d2af003c5150103c6050183c6250103c735012205518dc2066207d98e558d03c6550183c6450103c7650183c775012206558e4207e2075d8f598e0216518d2aec03c5950003c6850083c6a50003c7b5002205518dc2066207d98e558d03c6d50083c6c50003c7e50083c7f5002206558e4207e2075d8f598e0216518d2ae803c5150003c6050083c6250003c735002205518dc2066207d98e558d03c6550083c6450003c7650083c575002206558e4207e205d98dd18d82154d8d2ae413050002854597000000e780a09d630505422a8413060002814597100000e780e0d01145854597000000e780a09b63080540aa84a301050023010500a30005002300050013050002930b0002814597f0ffffe78060092a8bae8a2c001306000297100000e78060d9228597000000e780e09713054a0063634537814597f0ffffe7808006aae2aee682ea2320412dd00588028c0597f0ffffe780e0ee338649018802ce8597f0ffffe780e0ed166ab6695664268597000000e7804093dae2d6e6deead2eecef2a2f68545130514032308b116636a8530814597f0ffffe780c000aae4aee882ec0d4597d0ffffe780007f2330a12c2334b12c2338012c99c1814511a8880597e0ffffe780e08c8335012d0335012c8e052e95c1450ce18335012dd6698505138409012338b12c6362342d0335812c6399a500880597e0ffffe78080898335012d033a012c13953500529500e19384150005042338912c630f04280335812c639ca4008805a68597e0ffffe78060868334012d033a012c939a340033055a0100e136752295636d85262ad47010a8002c1097f0ffffe780c0de033b812c7d556384a4026410a10a52850c61130485002ed4a8002c10268697f0ffffe78060dce11a2285e3930afe63070b00528597000000e78060819665801a33863501a80097f0ffffe780e0d913061117a800a28597f0ffffe780e0d8f66536762e96a80097f0ffffe780e0d7a669c66a3665666a11c5166597f0ffffe780007d167511c5766597f0ffffe780207c82e002fc02f802f40403c802801a1306c002814597100000e78060ae130680132685814597100000e78060ad1775ffff930515cb4146228597100000e78000b9370501011b0505022320a114233c012a88051306800f814597100000e78020aa88058c0297b0ffffe78000b6a8008c051306800f97100000e78040b5a800ce85528697b0ffffe780c0bd8802ac001306800f97100000e78060b3880513060004814597100000e78080a5033581229305000263eaa50a5a655de5033501229a653386a50032e3ba66b335b600b6952ee78345012399c1fd552eeffd55130610082eeb637dc5121306000800136309c500098e2295814597100000e78040a088028402a28597b0ffffe78060c321459305312c9060a38ec5fe93568600238fd5fe93560601a38fd5fe935686012380d50093560602a380d500935686022381d50093560603a381d50061922382c5007d15a104a1055dfd0336812228108c0597100000e780a0a62c10130600024a8597100000e780a0a563870a004e8597f0ffffe780e0638330813f0334013f8334813e0339013e8339813d033a013d833a813c033b013c833b813b1301014082801775ffff1305e58825a01775ffff1305458839a81775ffff1305a58711a81775ffff1305058729a01775ffff13056586f14597e0ffffe780a02900001775ffff130525d89775ffff9386a5da9305b002900297e0ffffe780a04200001305000211a0114597f0ffffe780005c00009305000897f0ffffe780e09f0000697106f622f226ee4aea4ee652e2d6fddaf9def5e2f1e6ed2e8a2a89014481490d45aae082e49304110501163335c00093b51500b36ab500130b1108894b7d5c88088c0097f0ffffe780e056034501056309751f6301051003c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8d2ae903c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8d2ae503c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8d2ae103c5140083c5040003c6240083c6340022054d8d4206e206558e518d83c5540003c6440083c6640003c77400a205d18dc2066207d98ed58d82154d8daafc63890a00dda002e902e502e182fc639e0a0ca81813060002d28597100000e780c0c5012579e1639a091628110d46a28597e0ffffe780e0852a7559c96a75ca752a76aae9aee5b2e1a8188c0197f0ffffe78020320305eb008305db000346cb00e6792303a10aa205d18d2312b10a03459b0083458b000346ab008306bb0022054d8d4206e206558e518d2ad103451b0083450b0003462b0083463b0022054d8d4206e20683455b00558e518d03464b00a20583466b0003477b00d18d834c0108c2066207d98ed58d82154d8d2aed11a081496a658a550316410a8306610a2af82edc231ec102230fd102630e8409050401b5638609060305e1038315c1036256c2762307a1022316b10232d436f0130511010c103d4697000000e78080734ee423089101a8182c00054697f0ffffe78060eb667535c92a658a656676aaf0aeecb2e8880897f0ffffe78080012334a9004e8597f0ffffe78000b7014531a01305a005a300a90005452300a900b2701274f2645269b269126aee7a4e7bae7b0e7cee6c556182801775ffff1305c5a4f14597e0ffffe78000f700001775ffff130585ac9305b002edb71775ffff1305a5a49765ffff9386a52f9305b002900897e0ffffe780200f0000717106f522f126ed2a8432e402ec02e802fc02f8a303010232f4aee02800aae40808aae813057102aaec28109305710297f0ffffe780c02d058901e9034571020dc9a300a40005450da888102c101306800397000000e7804063f954ca65881097f0ffffe780c02a058969d991ccfd14f5b7c26562660ce810ec2300a400aa700a74ea644d61828097a0ffffe780c02d00004d7186e6a2e226fe4afa4ef652f256ee5aea5ee662e2e6fdeaf9eef5b2842e8a2ae0014c814d8149814b1304110cfd5a3d4d32e82ee48801e285268697d0ffffe780c04f0345010c631e052863045c3103459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8d2ae90345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8d2ae503459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8d2ae10345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8daafca81813060002d28597100000e780c08c0125631305188801e285268697d0ffffe780004d0e6b630d0b1ece6c2e65637f9d15aaeceef04145814597e0ffffe7800076aa84ae8b4146da8597000000e780204683c5840083c9940003caa40083cdb40003c6c40003cdd40083c7e40083caf40003c3040003c7140003ce240083c6340003c8440083c3540083c8640083c2740063870b04268542f4c68496e01a896af01e8d52ec728a6ef8b68dcee4ba89b2e856fcbe8aae8b97f0ffffe78060fede85d687e27a46664e87a669ee86c27d528e626aea83027d4a838662a68822780675631f0514a20933e5b900420ae20db3e54d014d8d220db365cd0013960701e20a33e6ca00d18d821533e9a500131587003365650093150e0113968601d18d4d8d93958300b3e505011396080193968201558ed18d82154d8daaf093840cff130a0b012685814597e0ffffe7802065aa8cae8bd285268697000000e7804035e6e1dee5a6e928118c0197f0ffffe78020e60c1988618c65814baa7daaf4aef88549c264226afd5a3d4d666511c55a8597f0ffffe780e0f0050c91bb2e6586765de533e5790111cd638c0d024675a675026608f20cee14e2233426012338b6013da01305500382652380a50023b80500638f0d006e8597e0ffffe780a07401a81305200382652380a50023b80500b6601664f2745279b279127af26a526bb26b126cee7c4e7dae7d716182801765ffff13054562f14597e0ffffe78080b400001765ffff130505639765ffff938685679305b002301197e0ffffe78080cd00001765ffff1305b56a93059002e9b797e0ffffe780c0cd0000757106e522e1a6fccaf8cef4d2f02a89814432e402e81304910181153335b00093351900b369b500094a28082c0097f0ffffe780a0e30345810165d9630c451303459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8daaec0345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8daae803459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8daae40345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8daae0e39909ee880013060002ca8597000000e78080530125e31e05ec93f4f40f850413f5f40fe30795ec1765ffff13058547f14597e0ffffe780c09900002685aa600a64e6744679a679067a4961828071c693f7f50f2300f5003307c500a30ff7fe894663fcc60aa300f5002301f500230ff7fea30ef7fe994663f1c60aa301f500230ef7fea14663fac60893f5f50f9b9785003307a0400d8bad9f198e9b950701ad9f2a97719a1cc3b305c70023aef5fe63f5c6065cc31cc723aaf5fe23acf5fee14663fcc604137847005cc71ccb5ccb1ccf6108939807029396070293d8080223a2f5fe23a4f5fe23a6f5fe23a8f5fe33060641fd474297c69663f0c7020116937706fe93870702ba9714e314e714eb14ef13070702e31af7fe8280397122fc26f84af44ef052ec56e85ae45ee093f735006387074069c2aa8719a06303062a83c60500850513f735002380d7007d1685076df793f637003e87cdea3d48637dc804930806ff6378180133e8b700137878006304083093d84800138f1800120f2e9f2e87be86832e0700032e4700032387000328c70023a0d60123a2c60123a4660023a606014107c106e31eeffc85089208c695c6973d8a137886001377460093762600058a630c080083a8050003a84500a107a10523ac17ff23ae07ff11c798419107910523aee7fe6391061e09c603c705002380e7006274c27422798279626ac26a226b826b216182807d476379c70a094883c805009841638806290d486386061d9306c6fe03c3150003c8250093f306ff13843700938435009382330123801701a38067002381070113d94600ae92a687a28803a8170083a5570083a697001b53870103a7d7009b1f88001b9f85009b9e86001b5888019bd585019bd686011b1e87003363f3013368e801b3e5d501b3e6c60123a0680023a2080123a4b80023a6d800c107c108e39657fa9307190092073516b385f40033067640a29793780601137886009376460013772600058a6384080883cb050003cb150083ca250003ca350083c9450003c9550083c4650003c4750083c3850083c2950083cfa50003cfb50083cec50003ced50003c3e50083c8f50023807701a380670123815701a381470123823701a382270123839700a383870023847700a38457002385f701a385e7012386d701a386c70123876700a3871701c105c1076304080483c2050083cf150003cf250083ce350003ce450003c3550083c8650003c8750023805700a380f7012381e701a381d7012382c701a382670023831701a3830701a105a1079dc203c3050083c8150003c8250083c6350023806700a380170123810701a381d70091059107e30307e283c6050003c715008907238fd7fea38fe7fe890539b513f73700e31d07ec39b59306c6fe93f306ff1384170093841500938213012380170113d94600ae92a687a28803a8370083a5770083a6b7001b53870003a7f7009b1f88011b9f85019b9e86011b5888009bd585009bd686001b1e87013363f3013368e801b3e5d501b3e6c60123a0680023a2080123a4b80023a6d800c107c108e39657fa9307190092073d16b385f40033067640a297a1b593d84800938e18002e88033e88000333080085062334c7012330670041084107e3e5d6ff85089208c695c6973d8a01bb9306c6fe03c8150093f306ff13842700938425009382230123801701a380070113d94600ae92a687a28803a8270083a5670083a6a7001b53070103a7e7009b1f08011b9f05019b9e06011b5808019bd505019bd606011b1e07013363f3013368e801b3e5d501b3e6c60123a0680023a2080123a4b80023a6d800c107c108e39657fa9307190092073916b385f40033067640a29749b3aa8709b919ca0347050083c705007d166317f700050585057df6014582800345050083c705001d9d8280aa862e87b287630db50cb388c5403308c040b388a84006082e832a8e6372181b3346b5001d8a637fb50a63010612cdcb1386f7ff9d4563f8c51813061700b305c54093b5750093c5150093f5f50f638a0516b365e5009d896395051693f587ffba95033603002103210e233ccefee39a65fe13f687ff13f57700aa87b385c600329739cd0345070005462380a5006389c704034517000946a380a5006382c704034527000d462381a500638bc702034537001146a381a5006384c7020345470015462382a500638dc700034557001946a382a5006386c700834767002383f5003685828029ea3306f5001d8a65ca1386f7fffdd7b307c5007d5821a07d16e30106ffb305c70003c5050093f57700fd17a380a700e5f59d4763fac70ab2871d48e117b305f7008861b385f60088e1e369f8fe93777600cdd7fd173306f700834506003386f6002300b600f5b71376750041ca9385f7ffc9d72a867d5821a0fd15e38005f903450700050693777600a30fa6fe0507edf79d4763fcb704938885ff93f888ffa10833051601ba8703b807002106a107233c06ffe31aa6fe469793f77500130617008ddfba9711a005060347f6ff0505a30fe5fee31af6fe36858280cdba3685d5b713061700f9bfb287a5b73285ae8713061700e1f919b73e8625bf2a86be8549bfd182e6ad7f520e5108c9bcf367e6096a1f6c3e2b8c68059b3ba7ca8485ae67bb6bbd41fbabd9831f2bf894fe72f36e3c79217e1319cde05bf1361d5f3af54fa54b598638d6c56d340101010101010101ff00ff00ff00ff00fffefefefefefefe80808080808080800a0a0a0a0a0a0a0a0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000018cd0900000000000010000000000000040000000000000018bd01000000000000100800000000004000000000000000010000000000000060090100000000000000000000000000011101250e1305030e10171b0eb44219110155170000023901030e0000032e001101120640186e0e030e3a0b3b053f198701190000042e00110112064018030e3a0b3b05360b3f198701190000052e006e0e030e3a0b3b05200b0000062e001101120640186e0e030e3a0b3b050000072e006e0e030e3a0b3b0b200b0000082e011101120640186e0e030e3a0b3b0b360b0000091d00311311011206580b590b570b00000a1d0031135517580b590b570b00000b1d00311311011206580b5905570b00000c1d0031135517580b5905570b00000d2e006e0e030e3a0b3b0b3f19200b00000e2e011101120640186e0e030e3a0b3b0b3f1900000f1d0131135517580b590b570b0000101d01311311011206580b590b570b0000111d01311311011206580b5905570b0000121d0131135517580b5905570b0000132e006e0e030e3a0b3b053f19200b0000142e011101120640186e0e030e3a0b3b05360b3f190000152e011101120640186e0e030e3a0b3b053f190000162e0111011206401831130000172e0011011206401831130000182e001101120640186e0e030e3a0b3b0b0000192e011101120640186e0e030e3a0b3b0b00001a2e011101120640186e0e030e3a0b3b0500001b2e011101120640186e0e030e3a0b3b05360b3f1987011900001c2e001101120640186e0e030e3a0b3b0b3f1987011900001d2e006e0e030e3a0b3b0b870119200b00001e2e001101120640186e0e030e3a0b3b0b360b3f198701190000007000000004000000000008016f2900001c001143000000000000051200000000000000000000700e0000021e2d00000200000000039a420100000000000e0000000152c44b000078350000010b0200021e2d000002463c000004a8420100000000000e00000001521d0e0000028e010300000000c722000004000000000008016f2900001c00f915000088000000051200000000000000000000a00e000002da180000021f050000057d0c00002f16000002f90501067877010000000000020000000152f03200002b0c000002eb01025c3c000002ab30000005fa350000712300000593030105fa350000712300000593030105fa350000712300000593030105fa350000712300000593030105fa35000071230000059303010594280000c52100000593030105e52a00001946000005930301056b380000833700000593030105c50b0000f90300000536050105fa3500007123000005930301000002ad0c000002ab300000055f3f00007123000007010401055f3f00007123000007010401055f3f00007123000007010401055f3f00007123000007010401055f3f0000712300000701040105c43000002c17000007010401054d0b0000e934000007010401000005a6000000c14600000273040105d71200000841000002730401056c4500002b050000024905010506080000cc000000024905010505280000f9030000026106010002a7300000023512000002a431000007454800004e27000003d00100022c3e0000071013000010460000038e0107403b0000a730000003890107403b0000a73000000389010000029c48000002632e0000087a770100000000004201000001529b1500008a35000004d3030965000000ea770100000000000200000004f1360adc1800000000000004f1150972000000fc770100000000000200000004f2360ae91800004000000004f215097f00000044780100000000000200000004fd360af61800007000000004fd1509f300000052780100000000000200000004fd470b000100006c78010000000000020000000403011e0b8c0000007e7801000000000002000000040701360c03190000a0000000040701150b0d0100008c7801000000000002000000040701470b1a0100009a7801000000000006000000040f0133000002a30b000007412b0000713b000004430107be2d0000482900000443010002242900000ddb130000b11b000004870100023c4400000d0d470000ce380000042a010002501400000e4880010000000000700000000152032e0000a7300000049a0fd902000020090000049b1110521a00004e8001000000000008000000044e1d11bd1900004e800100000000000800000019f8020909410100004e80010000000000080000001bef5000000af70200005009000004511c09d01e000060800100000000000400000004511609090300006e80010000000000080000000451280f952100008009000004651412071b0000b0090000225901090af41a0000e0090000171209000000000002650700000d87320000b11b000004870100026f0700000ed8860100000000007000000001521f030000a7300000049a0fe5020000800d0000049b1110a61a0000de8601000000000008000000044e1d11bd190000de860100000000000800000019f802090941010000de86010000000000080000001bef5000000ae2030000b00d000004511c09dd1e0000f086010000000000040000000451160909030000fe86010000000000080000000451280fa2210000e00d000004651412131b0000100e0000225901090af41a0000400e0000171209000000000000021f4a000013370a00006c0a000008bd0601137f030000672e000008f606011311490000f44000000810070105b90c000023050000086e050114bc78010000000000e4010000015289020000e031000008de04030bbc040000da780100000000000c00000008e504130bc9040000f6780100000000000400000008ea04190bd6040000327901000000000002000000080a051a12e3040000d00000000817052411c31c00001a7a010000000000040000000880051211b01c00001a7a010000000000040000000ec702090bfc1e00001a7a010000000000020000000e6d020c000000127511000010010000081a051112d01c0000400100000894041212b01c0000700100000ec702090cfc1e0000a00100000e6d020c00000012ac1e0000d0010000080b05200b50010000ac7901000000000006000000139403160b6a010000c07901000000000004000000139503090012b91e000000020000080c05210b5d010000b27901000000000004000000139403160b77010000c47901000000000004000000139503090011e3040000de790100000000001a000000080e052411c31c0000e479010000000000040000000880051211b01c0000e479010000000000040000000ec702090bfc1e0000e479010000000000040000000e6d020c00000011681d000008790100000000001c00000008eb041610031d000008790100000000001c00000012310910f71c000008790100000000001c000000112009105b1c000008790100000000001c00000011874c10ce1b000008790100000000001c00000010533111011c000008790100000000001c0000000a940d0910311c000008790100000000001c0000000c321110c11b000008790100000000001c0000000f7c091220190000300200000ab0091d1062190000147901000000000002000000092b350927010000147901000000000002000000095352000012431c0000800200000ab1091510711c00001679010000000000080000000f541c10141d000016790100000000000800000010501609bf1d000016790100000000000800000011871f000009121c00002079010000000000020000000f54150000000000000000000015f67a010000000000780300000152c0470000f92d0000083c0512701f0000b0020000083e05170c631f0000e00200001483020f00111a1e0000247b0100000000000400000008470525110d1e0000247b010000000000040000001641033311d0190000247b0100000000000400000016080327116e190000247b0100000000000400000019e502090999000000247b010000000000040000001b62500000000011e81b0000287b010000000000da0000000847052311db1b0000287b0100000000006e0000000a8b010912861d0000100300000a5801100f741d000040030000128c190fcb1d000070030000122c1209201900004c7b010000000000040000000b260e09e31d0000647b010000000000040000000b321209ef1d0000707b0100000000000a0000000b391309fb1d0000867b0100000000000a0000000b412509d71d0000607b010000000000040000000b2e1000000011dd1c0000487b010000000000040000000a57011211b01c0000487b010000000000040000000ec702090bfc1e0000487b010000000000020000000e6d020c00000011861d0000b47b0100000000004e0000000a8c010910741d0000b47b0100000000004a000000128c1910cb1d0000b47b0100000000004a000000122c120920190000b47b010000000000040000000b260e09fb1d0000ec7b0100000000000c0000000b412509ef1d0000e07b010000000000040000000b391309e31d0000dc7b010000000000040000000b32120000000012331e0000a0030000084c051312581e0000d003000016b9010911271e0000027c010000000000120000001814010c10dd190000087c0100000000000400000016dc1f0bbe1a0000087c01000000000004000000195a010f000000000c7d1f000000040000084c051c11681d0000367c010000000000720100000859052310031d0000367c0100000000007201000012310910f71c00003c7c0100000000001e000000112009105b1c00003c7c0100000000001e00000011874c10ce1b00003c7c0100000000001e00000010533111011c00003c7c0100000000001e0000000a940d0910311c00003c7c0100000000001e0000000c321110c11b00003c7c0100000000001e0000000f7c091220190000300400000ab0091d1062190000487c01000000000002000000092b350927010000487c01000000000002000000095352000012431c0000800400000ab1091510711c00004a7c010000000000080000000f541c10141d00004a7c0100000000000800000010501609bf1d00004a7c0100000000000800000011871f000009121c0000547c010000000000020000000f54150000000000000010211d00005a7c0100000000004e01000011220910ea1900005a7c01000000000014000000113a270b840100005a7c0100000000000600000019d60d1f11041a0000607c0100000000000800000019da0d200bf7190000607c0100000000000800000019460617000b111a0000687c0100000000000600000019db0d240010f71c00006e7c0100000000001a000000114715105b1c00006e7c0100000000001a00000011874c10ce1b00006e7c0100000000001a00000010533111011c00006e7c0100000000001a0000000a940d0910311c00006e7c0100000000001a0000000c321110c11b00006e7c0100000000001a0000000f7c091220190000b00400000ab0091d1062190000787c01000000000002000000092b350927010000787c01000000000002000000095352000012431c0000000500000ab1091510711c00007a7c010000000000080000000f541c10141d00007a7c0100000000000800000010501609bf1d00007a7c0100000000000800000011871f000009121c0000847c010000000000020000000f54150000000000000010f71c00008a7c0100000000001c000000114735105b1c00008a7c0100000000001c00000011874c10ce1b00008a7c0100000000001c00000010533111011c00008a7c0100000000001c0000000a940d0910311c00008a7c0100000000001c0000000c321110c11b00008a7c0100000000001c0000000f7c091220190000300500000ab0091d1062190000967c01000000000002000000092b350927010000967c01000000000002000000095352000012431c0000800500000ab1091510711c0000987c010000000000080000000f541c10141d0000987c0100000000000800000010501609bf1d0000987c0100000000000800000011871f000009121c0000a27c010000000000020000000f541500000000000000102d1d0000dc7c01000000000012000000115a1209e91f0000e87c01000000000004000000117f0e0010ab1900000a7d01000000000006000000115019102b1a00000a7d010000000000060000001b1a0e117a1900000a7d0100000000000600000019e5020909a60000000a7d010000000000060000001b62500000000a2c190000b00500001150190a391d0000f005000011541b0f381900006006000011631a10861900007c7d01000000000002000000092b3509340100007c7d01000000000002000000095352000009451d00007e7d0100000000000c00000011641b10511d0000947d0100000000001200000011661609f61f0000a07d01000000000004000000117f0e00091e1a0000067d01000000000004000000114f2c1098190000f27c01000000000010000000114a12114b1f0000fe7c010000000000040000001bcb051b113d1f0000fe7c010000000000040000000d7e04080b2b1f0000fe7c010000000000040000000d2e030900000000000012e3040000b00600000863052811c31c0000047e010000000000040000000880051211b01c0000047e010000000000040000000ec702090bfc1e0000047e010000000000020000000e6d020c0000001175110000307e010000000000260000000865051512d01c0000f00600000894041212b01c0000200700000ec702090cfc1e0000500700000e6d020c000000000d3c380000ae2d000008f2011337170000372b000008f4050113263100001729000008430701051a270000431c0000089c0401167a850100000000009800000001526211000011f916000086850100000000001800000008e6071b0b6510000086850100000000000c0000001f1701120011c1160000ac850100000000005800000008e807091169210000b6850100000000004a0000001f65012711b5150000b885010000000000480000002027051611c9150000cc85010000000000060000001f66013c0bc9040000cc85010000000000060000001f700109000b65100000d485010000000000140000001f6701150b65100000ea85010000000000160000001f69011100000000131f0700005723000008e5070100021e1a000005f8160000fb2e0000089304010002012f000002e031000006a07a010000000000560000000152cf490000d819000008f304000005fa0800008b49000008640401051b0f00001f09000008790401157c7e0100000000007e010000015245390000fb2e00000838040c591000008007000008390419128b1c0000b0070000084d041d0a44190000e00700001d2f110012a9110000100800000856041a11b6110000047f01000000000018000000086b04150bb30100000a7f010000000000120000000881042c0011b61100002a7f01000000000018000000086c04190bb3010000307f010000000000120000000881042c0011381a00004a7f010000000000040000000873041f11ca1a00004a7f010000000000040000001996011a09b30000004a7f0100000000000400000017ee1c00000bbf0100004e7f010000000000080000000876040b0012971c000040080000083f041d0a50190000700800001d2f11000bcb0100009c7f0100000000000a0000000846041512451a0000a0080000085d042612d61a0000e0080000195a010f10e21a0000ca7f0100000000000400000017d93609c0000000ca7f0100000000000400000017ee1c0000000002f101000007d53c0000bd3800001f550102ec3700000eb880010000000000bc010000015292350000372b00001f1f0fab1d0000100a00001f201212981d0000400a0000123f050911971e00003e81010000000000d40000001272020f116c1a0000488101000000000008000000249e01320b251b0000488101000000000008000000195a010900116f1b00005081010000000000ac00000024a20122097b1b000056810100000000001a000000252c1010871b000070810100000000008c000000252f0510cd00000070810100000000000c0000002552160b8401000070810100000000000c0000000540051600109f1b0000b6810100000000000a000000256a160910200000b681010000000000020000002514070010931b0000a0810100000000000a0000002569160903200000a081010000000000020000002514070009da00000094810100000000000400000025651b097b1b0000e88101000000000014000000257716097b1b0000c88101000000000012000000255a1e000011791a000008820100000000000200000024b701430b251b0000088201000000000002000000195a010900111c1f00000a820100000000000400000024b8011c115c1b00000a82010000000000040000000da9050d093e1b00000a8201000000000004000000231a0900000000000f401e0000700a00001f252712841e0000a00a0000165f040d12711e0000d00a000024450229125f1a0000000b000024de0309110f1f00001a810100000000000a0000001909091311501b00001a810100000000000a0000000da9050d093e1b00001a810100000000000a000000231a09000000000000000002623d000002f644000005920400004e2700001f3501010002d119000005fc2200004e2700001f6501010000023d290000058f490000ae4600001f6f0101155a84010000000000200100000152bd090000f64400001f3401125c210000b00b00001f35012311a21500007e84010000000000de0000002027051612c9150000e00b00001f3601100cc9040000100c00001f700109000b65100000a684010000000000160000001f3801150c65100000400c00001f4101110b7c210000dc84010000000000020000001f41011112d4160000700c00001f3c01220f7f100000b00c00001f1a0911eb160000fc840100000000000a00000008a30412098a1f0000fc840100000000000a0000001f1a260000000b651000004885010000000000120000001f3e011100000013bd1c0000d11900001f6301010002b547000007821c0000b92d00001f15010002f108000002b92d0000071f3500004e2700001f1a0100000569310000ec2200001f1301010002e82f0000167482010000000000b400000001526b17000010b922000082820100000000009600000008a41a11a72200008282010000000000960000002679022a0c9a220000300b000026b6060f00000017288301000000000038000000015277170000074d180000ee2f000008a30107c5440000994b000008bf010002ab3000001860830100000000000a0000000152ef4700002842000008c6196a83010000000000b6000000015253420000ee2f000008ca106b1700007883010000000000a200000008cb0910b92200007a830100000000009600000008a41a11a72200007a83010000000000960000002679022a0c9a220000700b000026b6060f000000001920840100000000003a000000015296370000994b000008ce097717000040840100000000001400000008cf090000027809000005b40f0000a730000008bb09010002210c00001a20860100000000001600000001525f300000ff0f000008d0080b3d18000020860100000000001600000008d0083e000000028c39000002164a0000029548000019747701000000000004000000015282090000fd4b000001fa10a101000074770100000000000400000001fa05093400000074770100000000000200000003d21e0000000000029039000005f909000068100000065f0a0105f909000068100000065f0a0105f909000068100000065f0a0105f909000068100000065f0a010002b131000002fa1c00000279230000077a33000056450000097c0107c63a0000c1010000097c01076b2a000027410000097c0107b34a00000b3e0000097c0107f91a0000b73c0000097c0100024c3600000712000000fd190000094b01072b2d0000514900001b5b0107f5310000d52100001b5b0107e52100005f340000094b010002a94a00000503370000274100001bc705010002ab30000007c20a0000b03a00001b190100029b0b000007731b0000dd4100001bd901000002ab30000005641100002a1a000019e4020105a91a0000f62700001956010105f1430000e246000019cb0d010585250000ac3d00001998060105b3050000c33d0000194206010543410000b008000019860d010534280000802800001916040105f53700009f3a000019e402010553190000ab110000198f01010597410000432f000019560101051f2600002809000019f7020105a90d0000ca17000019040901054c040000a919000019560101054c040000a919000019560101020f0700000312860100000000000e0000000152ab4200007a390000190b0d00051f2600002809000019f702010002b403000002ec370000074a050000ed31000017d7010775340000f028000017e30107400d0000d911000017d70107353e00001231000017e30100028d37000005fa0100003646000017ec01010002ab30000007542f00006c17000017110107542f00006c1700001711010002623d000005c3140000ed310000175f0101000002ec0c00000259490000075a140000983b00002352010002ab30000007b71b0000573d000023190107b71b0000573d0000231901000002b22d000007d8170000b22d000025290107a63b0000de3b00002534010d74470000341c000025470107760f0000a93e000025130107760f0000a93e0000251301000002fa1c000002242d000002b029000002494300000538120000842300000aaa090105663c0000ad3f00000a8f0d01058f360000f60000000a560101053a080000ba0e00000a8a0101000002801000000286100000075a2700009b3900000c310102b50c00000780400000901000000c35010000000002b846000002712e000002ec37000007752e0000ff1c00000f78010002304a0000075e4300001c1f00000f5401000002294a000002ec370000077907000078120000104d01020c000000025f4500000744160000590000001050010000000002ef1a000002f108000007fe050000db2500001d2e0107461300002c2200001d2e01000000022d08000002ec3700000593450000ca2000000e6c02010002cc46000005db200000274100000ec6020105db200000274100000ec6020105db200000274100000ec602010000000208000000020c0000000d760a0000e519000011860107270e000052430000111a0102e519000007be1e00004e270000118701000d790800004419000011260107d03d0000fd120000117a0107242a0000d201000011720107242a0000d201000011720107d03d0000fd120000117a010002fa1c000002ab30000007a04800000c00000012300107394a00001f01000012290100025949000007331a00001f010000128a010002cf2f00000570260000b00b0000126c020100020b42000005e22b0000dd2f0000123e0501000002b60a0000076b3d0000a53c00000b180107b9290000d63600000b240107dc0e0000f82900000b0b010770210000b22100000b11010770210000b22100000b11010770210000b22100000b11010002ab3000000551360000f73300001607030105b0270000d54600001640030107f60c0000082a000016d30105fd3300003934000016b80101050a040000473d0000165b04010002242d000002bb300000052401000046050000181301010000025f4700000224290000052d4b00006747000024dd03010002cc46000005be26000067470000244102010002ab30000005642c00003a320000249b0101000000026845000005673a0000101a0000138f030105b73100005b0e0000138f0301027c2b00000244140000056e4400000347000021e80101056e4400000347000021e8010100000002ec0c000002f00c000002ec00000005df180000f43300000d5305010002e322000005d43800002e2900000da8050105d43800002e2900000da80501000005464400000a2f00000d930401027f3700000562490000192a00000d2a03010005cc080000192a00000d7d040100023308000002b4300000057d0e0000370500001456020105b4430000903a00001482020105ba0300003341000014bb03010591060000f50d000014120601001b2c800100000000000e00000001522c3f00006c390000148b070311492000002e800100000000000c000000148c0705093d2000002e800100000000000c0000001c8605000000029c480000023c44000005662d0000f64600001ae4040105662d0000f64600001ae4040105664600008c4b00001acd040105664600008c4b00001acd0401000002e62800001c6e7e0100000000000e0000000152cc150000fd2d00001c6e1d113d0000e31100001c95011d450f00005f3100001c85011e3a800100000000000e000000015224300000154200001c50030002a4190000021526000015fa7f010000000000120000000152fc440000a73000001ebb021172100000fa7f010000000000120000001ebc021b1137130000fa7f01000000000012000000084407090965100000fa7f010000000000120000001f5912000000000230320000150c80010000000000120000000152c2020000a73000001ed60211721000000c80010000000000120000001ed7021b11371300000c80010000000000120000000844070909651000000c80010000000000120000001f5912000000000002d4130000031e800100000000000e0000000152ec040000f711000020720602ae4700000545320000801800002025050105cd060000eb3b00002025050100021a30000005bc3e00005b090000209b07010000026a26000002c01700000563220000892b0000225801010563220000892b00002258010100021a3000000e3686010000000000a2000000015207100000a730000022830f62110000f00c000022830a12f9160000200d000008e6071b0c65100000500d00001f1701120011c116000074860100000000005800000008e8070911692100007e860100000000004a0000001f65012711b51500008086010000000000480000002027051611c91500009486010000000000060000001f66013c0bc90400009486010000000000060000001f700109000b651000009c86010000000000140000001f6701150b65100000b286010000000000160000001f69011100000000000000028c060000021735000005db2c0000091800002699060105121800000e2d000026b5060102ab300000054c150000b94400002677020100000000003c0000000200000000000800ffffffff9a420100000000000e00000000000000a8420100000000000e0000000000000000000000000000000000000000000000bc0100000200740000000800ffffffff74770100000000000400000000000000787701000000000002000000000000007a770100000000004201000000000000bc78010000000000e401000000000000a07a0100000000005600000000000000f67a01000000000078030000000000006e7e0100000000000e000000000000007c7e0100000000007e01000000000000fa7f01000000000012000000000000000c8001000000000012000000000000001e800100000000000e000000000000002c800100000000000e000000000000003a800100000000000e0000000000000048800100000000007000000000000000b880010000000000bc010000000000007482010000000000b4000000000000002883010000000000380000000000000060830100000000000a000000000000006a83010000000000b60000000000000020840100000000003a000000000000005a8401000000000020010000000000007a85010000000000980000000000000012860100000000000e00000000000000208601000000000016000000000000003686010000000000a200000000000000d886010000000000700000000000000000000000000000000000000000000000ec77010000000000f077010000000000f477010000000000fc7701000000000008780100000000000c7801000000000000000000000000000000000000000000fe7701000000000006780100000000000c780100000000001478010000000000000000000000000000000000000000004678010000000000527801000000000054780100000000005e780100000000000000000000000000000000000000000080780100000000008c780100000000008e7801000000000096780100000000000000000000000000000000000000000036790100000000003c7901000000000040790100000000004679010000000000fa790100000000002a7a010000000000000000000000000000000000000000005a7a0100000000007a7a0100000000009a7a010000000000a07a01000000000000000000000000000000000000000000627a0100000000006a7a0100000000009a7a010000000000a07a01000000000000000000000000000000000000000000627a0100000000006a7a0100000000009a7a010000000000a07a01000000000000000000000000000000000000000000627a0100000000006a7a0100000000009a7a010000000000a07a01000000000000000000000000000000000000000000ac79010000000000b279010000000000c079010000000000c47901000000000000000000000000000000000000000000b279010000000000b679010000000000c479010000000000c8790100000000000000000000000000000000000000000008790100000000000c79010000000000147901000000000016790100000000001e790100000000002079010000000000227901000000000024790100000000000000000000000000000000000000000016790100000000001e790100000000002079010000000000227901000000000000000000000000000000000000000000f87a0100000000000e7b010000000000107b010000000000187b01000000000000000000000000000000000000000000f87a0100000000000e7b010000000000107b010000000000187b010000000000000000000000000000000000000000003a7b010000000000447b0100000000004c7b010000000000967b010000000000000000000000000000000000000000003a7b0100000000003e7b0100000000004c7b010000000000927b010000000000000000000000000000000000000000003a7b0100000000003e7b0100000000004c7b010000000000927b01000000000000000000000000000000000000000000027c010000000000187c0100000000001e7c010000000000227c01000000000000000000000000000000000000000000027c010000000000187c0100000000001e7c010000000000227c010000000000000000000000000000000000000000001a7c0100000000001e7c010000000000247c010000000000267c010000000000000000000000000000000000000000003c7c010000000000407c010000000000487c0100000000004a7c010000000000527c010000000000547c010000000000567c0100000000005a7c010000000000000000000000000000000000000000004a7c010000000000527c010000000000547c010000000000567c010000000000000000000000000000000000000000006e7c010000000000727c010000000000787c0100000000007a7c010000000000827c010000000000847c010000000000867c010000000000887c010000000000000000000000000000000000000000007a7c010000000000827c010000000000847c010000000000867c010000000000000000000000000000000000000000008a7c0100000000008c7c010000000000967c010000000000987c010000000000a07c010000000000a27c010000000000a47c010000000000a67c01000000000000000000000000000000000000000000987c010000000000a07c010000000000a27c010000000000a47c01000000000000000000000000000000000000000000107d010000000000127d010000000000567d0100000000005a7d0100000000005c7d010000000000627d010000000000000000000000000000000000000000001a7d010000000000227d010000000000247d010000000000287d0100000000002a7d010000000000307d010000000000327d010000000000427d010000000000447d010000000000467d0100000000004a7d010000000000567d01000000000000000000000000000000000000000000627d0100000000007a7d0100000000007c7d0100000000007e7d0100000000008a7d0100000000008c7d0100000000008e7d010000000000927d01000000000000000000000000000000000000000000ac7d010000000000b27d010000000000b67d010000000000bc7d010000000000e27d010000000000147e01000000000000000000000000000000000000000000387e010000000000407e010000000000527e010000000000567e01000000000000000000000000000000000000000000387e010000000000407e010000000000527e010000000000567e01000000000000000000000000000000000000000000387e0100000000003c7e010000000000527e010000000000567e01000000000000000000000000000000000000000000947e0100000000009c7e010000000000a07e010000000000a87e01000000000000000000000000000000000000000000ae7e010000000000d87e010000000000587f010000000000687f01000000000000000000000000000000000000000000ae7e010000000000d87e010000000000587f010000000000687f01000000000000000000000000000000000000000000ea7e010000000000f87e010000000000fc7e010000000000567f010000000000000000000000000000000000000000006c7f0100000000008a7f010000000000a87f010000000000b27f010000000000000000000000000000000000000000006c7f0100000000008a7f010000000000a87f010000000000b27f01000000000000000000000000000000000000000000b67f010000000000bc7f010000000000c27f010000000000c67f010000000000ca7f010000000000ce7f01000000000000000000000000000000000000000000b67f010000000000bc7f010000000000c27f010000000000c67f010000000000ca7f010000000000ce7f010000000000000000000000000000000000000000004e80010000000000a480010000000000aa80010000000000b880010000000000000000000000000000000000000000005e80010000000000608001000000000076800100000000007a800100000000000000000000000000000000000000000084800100000000008e80010000000000aa80010000000000b8800100000000000000000000000000000000000000000084800100000000008e80010000000000aa80010000000000b8800100000000000000000000000000000000000000000084800100000000008e80010000000000aa80010000000000b88001000000000000000000000000000000000000000000fe8001000000000016810100000000003681010000000000128201000000000000000000000000000000000000000000fe8001000000000016810100000000003681010000000000128201000000000000000000000000000000000000000000168101000000000024810100000000004282010000000000468201000000000000000000000000000000000000000000168101000000000024810100000000004282010000000000468201000000000000000000000000000000000000000000168101000000000024810100000000004282010000000000468201000000000000000000000000000000000000000000168101000000000024810100000000004282010000000000468201000000000000000000000000000000000000000000828201000000000086820100000000008e820100000000009482010000000000b082010000000000b682010000000000000000000000000000000000000000007a830100000000007e8301000000000086830100000000008c83010000000000a883010000000000ae8301000000000000000000000000000000000000000000708401000000000072840100000000007e840100000000005c8501000000000000000000000000000000000000000000828401000000000086840100000000008a840100000000008e8401000000000000000000000000000000000000000000828401000000000086840100000000008a840100000000008e8401000000000000000000000000000000000000000000cc84010000000000d684010000000000d884010000000000dc8401000000000000000000000000000000000000000000ea84010000000000ee84010000000000f48401000000000032850100000000003685010000000000408501000000000000000000000000000000000000000000ea84010000000000ee84010000000000f48401000000000032850100000000003685010000000000408501000000000000000000000000000000000000000000408601000000000042860100000000004486010000000000cc8601000000000000000000000000000000000000000000408601000000000042860100000000004486010000000000608601000000000000000000000000000000000000000000408601000000000042860100000000004486010000000000548601000000000000000000000000000000000000000000de8601000000000034870100000000003a87010000000000488701000000000000000000000000000000000000000000ee86010000000000f08601000000000006870100000000000a870100000000000000000000000000000000000000000014870100000000001e870100000000003a8701000000000048870100000000000000000000000000000000000000000014870100000000001e870100000000003a8701000000000048870100000000000000000000000000000000000000000014870100000000001e870100000000003a870100000000004887010000000000000000000000000000000000000000009a42010000000000a842010000000000a842010000000000b642010000000000000000000000000000000000000000007477010000000000787701000000000078770100000000007a770100000000007a77010000000000bc78010000000000bc78010000000000a07a010000000000a07a010000000000f67a010000000000f67a0100000000006e7e0100000000006e7e0100000000007c7e0100000000007c7e010000000000fa7f010000000000fa7f0100000000000c800100000000000c800100000000001e800100000000001e800100000000002c800100000000002c800100000000003a800100000000003a8001000000000048800100000000004880010000000000b880010000000000b8800100000000007482010000000000748201000000000028830100000000002883010000000000608301000000000060830100000000006a830100000000006a83010000000000208401000000000020840100000000005a840100000000005a840100000000007a850100000000007a85010000000000128601000000000012860100000000002086010000000000208601000000000036860100000000003686010000000000d886010000000000d8860100000000004887010000000000000000000000000000000000000000007261775f7665630073747200636f756e74005f5a4e34636f726535736c6963653469746572313349746572244c542454244754243134706f73745f696e635f73746172743137683231633736663939343638653065646545007b636c6f7375726523307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e005f5a4e34636f726533707472347265616431376831626239643039646638396234373532450077726974653c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e007b696d706c2335347d00616476616e63655f62793c636f72653a3a7374723a3a697465723a3a43686172496e64696365733e006e657874005f5a4e34636f726533737472367472616974733131305f244c5424696d706c2475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c5424737472244754242475323024666f722475323024636f72652e2e6f70732e2e72616e67652e2e52616e6765546f244c54247573697a652447542424475424336765743137683633326532303137643665353735396645006e6578743c5b7573697a653b20345d3e00636f6e7461696e735f6e6f6e5f636f6e74696e756174696f6e5f62797465006275696c64657273005f5a4e3131305f244c5424636f72652e2e6f70732e2e72616e67652e2e52616e676546726f6d244c54247573697a6524475424247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c54242475356224542475356424244754242447542435696e6465783137686163396536316662616530626263376145005f5a4e34636f726533666d7439466f726d617474657231327061645f696e74656772616c3137686238656639343965396131613633346545005f5a4e36335f244c5424636f72652e2e63656c6c2e2e426f72726f774d75744572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683636336332373865383138373636393045005f5a4e34636f726533666d74336e756d35335f244c5424696d706c2475323024636f72652e2e666d742e2e55707065724865782475323024666f7224753230246936342447542433666d743137683464336136353331313038303933376445005f5a4e34636f726533666d7439466f726d617474657239616c7465726e617465313768333537326537646636323036356664374500696e646578005f5a4e34636f7265366f7074696f6e31354f7074696f6e244c5424542447542439756e777261705f6f72313768343165333439646137383638346138334500616c69676e5f6f66667365743c75383e005f5a4e34636f72653373747232315f244c5424696d706c24753230247374722447542439656e64735f776974683137683139626662313333653233336465306145005f5a4e34636f726535736c69636532395f244c5424696d706c2475323024247535622454247535642424475424336765743137683233646638653962656438656665346645005f5a4e34636f726533666d74386275696c64657273313044656275675475706c65356669656c6432385f24753762242475376224636c6f73757265247537642424753764243137686363643963626231656235626135633645005f5a4e34636f726536726573756c743133756e777261705f6661696c65643137683030653934303161326339653536633045007074720070616464696e670077726974653c636861723e0069735f736f6d653c7573697a653e00676574005f5a4e37355f244c54247573697a65247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c542424753562245424753564242447542424475424336765743137683362336666656535366439303731313345005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243873706c69745f61743137683461343239666364306233623563343945005f5a4e3131305f244c5424636f72652e2e697465722e2e61646170746572732e2e656e756d65726174652e2e456e756d6572617465244c54244924475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e65787431376831623734616564656639323065303665450063686172005f5a4e34636f7265366f7074696f6e31354f7074696f6e244c5424542447542436696e736572743137686265366237313331636461646331646245005f5a4e34636f726536726573756c743139526573756c74244c542454244324452447542438616e645f7468656e313768316532623263316238653933626561654500636f70795f66726f6d5f736c696365005f5a4e34636f726533666d7439466f726d6174746572323564656275675f7475706c655f6669656c64315f66696e6973683137683963326264643732306464613133376545007b696d706c2332397d007b696d706c2336357d005f5a4e3130385f244c5424636f72652e2e697465722e2e61646170746572732e2e66696c7465722e2e46696c746572244c5424492443245024475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722447542435636f756e743137683631323362313132363938303130326445005f5a4e34636f72653370747235777269746531376830336462313664353065636536366165450072616e6765006f7074696f6e005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f72336e74683137683635613666633036633265613031396645005f5a4e34636f72653373747235636f756e743134646f5f636f756e745f6368617273313768653066306166323562653730356463664500616c69676e5f746f5f6f6666736574733c75382c207573697a653e005f5a4e34636f726533636d70336d696e3137683961303232643031326665326338333745007b696d706c23317d005f5a4e34636f726533666d743372756e313768666639613633333362396633663061614500676574636f756e7400697465725f6d75743c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e006272616e63683c28292c20636f72653a3a666d743a3a4572726f723e007b696d706c2332357d005f5a4e34636f7265336f70733866756e6374696f6e36466e4f6e63653963616c6c5f6f6e63653137683331326365396462383432326365623645005f5a4e34636f726533666d74386275696c64657273313044656275675475706c65356669656c643137686134393061356537663734366534656245005f5a4e34636f72653130696e7472696e736963733139636f70795f6e6f6e6f7665726c617070696e673137683165326664363834393232323263326345005f5a4e34636f726533666d7439466f726d6174746572397369676e5f706c75733137683765363563323535316433616561343445007369676e5f706c7573005f5a4e34636f72653373747235636f756e743233636861725f636f756e745f67656e6572616c5f6361736531376864313333363866323830386530613030450076616c69646174696f6e73005f5a4e34636f726535736c696365346974657238375f244c5424696d706c2475323024636f72652e2e697465722e2e7472616974732e2e636f6c6c6563742e2e496e746f4974657261746f722475323024666f7224753230242452462424753562245424753564242447542439696e746f5f697465723137683765326332623733366531386264656545005f5a4e34636f726533707472376d75745f70747233315f244c5424696d706c2475323024244250246d75742475323024542447542433616464313768333939313037663564323335643062374500497465724d75740047656e657269635261646978006e6578745f696e636c75736976653c636861723e005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243132616c69676e5f6f66667365743137686265366661383332613635626436303545007b696d706c2335337d0064726f705f696e5f706c6163653c26636f72653a3a697465723a3a61646170746572733a3a636f706965643a3a436f706965643c636f72653a3a736c6963653a3a697465723a3a497465723c75383e3e3e005f5a4e34636f7265337074723133726561645f766f6c6174696c653137683034656338646164326362346562306245006d75745f7074720073756d005f5a4e34636f726533666d7439466f726d61747465723770616464696e67313768386664646163386139653836623737364500636d7000696d706c73005f5a4e34636f72653373747232315f244c5424696d706c247532302473747224475424313669735f636861725f626f756e646172793137683034353265303532643135616334353245005f5a4e37355f244c54247573697a65247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c542424753562245424753564242447542424475424336765743137686337356165633633323166633531643545005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542439656e64735f77697468313768383363653331633938643238356662364500696e736572743c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e005f5f72646c5f6f6f6d005f5a4e34636f72653373747235636f756e743131636f756e745f63686172733137683362393037393633646461313835376345007265706c6163653c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e005f5a4e34636f7265366f7074696f6e31354f7074696f6e244c542454244754243769735f736f6d653137686166353061376333383437653666373645006e74683c636f72653a3a7374723a3a697465723a3a43686172496e64696365733e005f5a4e34636f726533737472313176616c69646174696f6e733135757466385f66697273745f627974653137683962396637633933306431356335663945005f5a4e34636f726533666d7438676574636f756e743137683639663830313763343363306364653245005f5a4e34636f72653970616e69636b696e673970616e69635f7374723137683666303932373830653338346562353045005f5a4e34636f726535736c696365366d656d6368723138636f6e7461696e735f7a65726f5f627974653137686130353638656531383330306135373245005f5a4e34355f244c5424244c502424525024247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d74313768613430323766643039663261636331324500666d743c28293e005f5a4e36375f244c5424636f72652e2e61727261792e2e54727946726f6d536c6963654572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d74313768353264643636336235383463633535664500636f70795f6e6f6e6f7665726c617070696e673c75383e00616363756d007b696d706c2334387d007b636c6f7375726523307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542434697465723137686266616536663139613561623764656445006765745f756e636865636b65643c636f72653a3a666d743a3a72743a3a417267756d656e742c207573697a653e006765743c267374723e0070616e69635f646973706c61793c267374723e00756e777261705f6661696c6564002f72757374632f32663662633564323539653761623235646466646433336465353362383932373730323138393138007274005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f7234666f6c64313768623061333862663336373733633236364500636f756e743c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e005f5a4e34636f726533707472347265616431376831653634383335653639376533366630450073756d5f62797465735f696e5f7573697a65005f5a4e34636f726533666d7432727438417267756d656e743861735f7573697a653137686437613231613332353662616362386245005f5a4e3131305f244c5424636f72652e2e697465722e2e61646170746572732e2e656e756d65726174652e2e456e756d6572617465244c54244924475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e657874313768633030313137313163643937383139624500726573756c74005f5a4e37335f244c5424636f72652e2e666d742e2e6e756d2e2e4c6f776572486578247532302461732475323024636f72652e2e666d742e2e6e756d2e2e47656e657269635261646978244754243564696769743137686634306237613733623764393162653445004d61796265556e696e6974007b696d706c2336347d005f5a4e37335f244c54242475356224412475356424247532302461732475323024636f72652e2e736c6963652e2e636d702e2e536c6963655061727469616c4571244c542442244754242447542435657175616c3137686637383434376536346661643333376145005f5a4e3130365f244c5424636f72652e2e6f70732e2e72616e67652e2e52616e6765244c54247573697a6524475424247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c542424753562245424753564242447542424475424336765743137683761383664333261616263343034303345005f5a4e34636f72653463686172376d6574686f647332325f244c5424696d706c247532302463686172244754243131656e636f64655f757466383137683661333732316366346263313738623645005f5a4e34636f726533666d74336e756d33696d7037666d745f7536343137683238366534643532373433386334363745005f5a4e34636f72653970616e69636b696e673570616e69633137686437373538656430613265383739363145006c6962726172792f636f72652f7372632f6c69622e72732f402f636f72652e353431663036343835316338633866372d6367752e3000726561645f766f6c6174696c653c7573697a653e005f5a4e3130385f244c5424636f72652e2e697465722e2e61646170746572732e2e66696c7465722e2e46696c746572244c5424492443245024475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722447542435636f756e7438746f5f7573697a6532385f24753762242475376224636c6f73757265247537642424753764243137686532646263323632336436376436643345005f5a4e34636f726533666d743131506f737450616464696e673577726974653137683130373832303864313037663934393045006164643c7573697a653e005f5a4e34636f726533666d7439466f726d61747465723977726974655f737472313768353330393765363135313339346565644500696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e2c20636f72653a3a6f70733a3a72616e67653a3a52616e676546726f6d3c7573697a653e3e007b696d706c2331357d00656e64735f776974683c75383e005f5a4e34636f726535736c696365366d656d636872366d656d6368723137683838333063653264646237323666636245006c656e5f75746638005f5a4e34636f72653463686172376d6574686f64733135656e636f64655f757466385f7261773137686230336466376165346464366562316445005f5a4e34636f726533666d74355772697465313077726974655f63686172313768666466623438666364333637346132384500616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23347d3a3a6669656c643a3a7b636c6f737572655f656e7623307d3e00636f7265005f5a4e34636f726533636d7035696d706c7335375f244c5424696d706c2475323024636f72652e2e636d702e2e5061727469616c4f72642475323024666f7224753230247573697a6524475424326c74313768383563303932356636663163316566654500646f5f636f756e745f6368617273005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542431336765745f756e636865636b656431376838333832313033623533356331333034450063656c6c006765743c75382c20636f72653a3a6f70733a3a72616e67653a3a52616e67653c7573697a653e3e0066696e6973680077726974655f70726566697800636861725f636f756e745f67656e6572616c5f6361736500706f73745f696e635f73746172743c75383e007265706c6163653c636861723e00506f737450616464696e6700697465723c75383e005f5a4e38375f244c5424636f72652e2e7374722e2e697465722e2e43686172496e6469636573247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683862646365633661316137393933386345005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542433676574313768396431656137353833353464396166364500656e756d6572617465005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683563636236663439653430616432356245005f5a4e34636f726535736c69636534697465723136497465724d7574244c54245424475424336e65773137683131393134666634646337396132326545006469676974005f5a4e34636f726535736c69636533636d7038315f244c5424696d706c2475323024636f72652e2e636d702e2e5061727469616c4571244c54242475356224422475356424244754242475323024666f7224753230242475356224412475356424244754243265713137683331383339323064643563373930336445006d656d6368725f616c69676e656400777261705f6275663c636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23317d3a3a777261703a3a7b636c6f737572655f656e7623307d3e005f5a4e34636f726533666d74386275696c6465727331305061644164617074657234777261703137686630613261643433323636313138356545005f5a4e34636f726533666d74386275696c64657273313044656275675475706c653666696e6973683137683262326465366164386361323965353845006974657200666f6c643c7573697a652c20636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c207573697a652c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e005f5a4e34636f72653373747235636f756e743233636861725f636f756e745f67656e6572616c5f6361736532385f24753762242475376224636c6f73757265247537642424753764243137686238333838383631636166343538396545007b636c6f7375726523307d3c2675382c207573697a652c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e00737065635f6e6578743c7573697a653e005f5a4e34636f726534697465723572616e67653130315f244c5424696d706c2475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722475323024666f722475323024636f72652e2e6f70732e2e72616e67652e2e52616e6765244c5424412447542424475424346e6578743137683166316635393732633862353338396245005f5a4e34636f726533737472313176616c69646174696f6e733138757466385f6163635f636f6e745f62797465313768386431353839303565613233346333334500757466385f6163635f636f6e745f62797465006164643c5b7573697a653b20345d3e006e65773c5b7573697a653b20345d3e005f5a4e34636f726535736c6963653469746572313349746572244c542454244754243134706f73745f696e635f73746172743137686632323465323937613136633263656145006e6578743c636f72653a3a736c6963653a3a697465723a3a497465723c636f72653a3a666d743a3a72743a3a417267756d656e743e3e005f5a4e34636f726535617272617938355f244c5424696d706c2475323024636f72652e2e6f70732e2e696e6465782e2e496e646578244c542449244754242475323024666f722475323024247535622454247533622424753230244e24753564242447542435696e6465783137683663646534633833393961376530333445007b696d706c23397d0064656275675f7475706c655f6e6577005f5a4e34636f726533666d74386275696c64657273313044656275675475706c653666696e69736832385f24753762242475376224636c6f737572652475376424247537642431376861393666623161373161643166373535450064656275675f7475706c655f6669656c64315f66696e697368006164643c75383e007b696d706c233138317d00666f6c643c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a6d61703a3a6d61705f666f6c643a3a7b636c6f737572655f656e7623307d3c2675382c207573697a652c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e3e005f5a4e34636f726535736c69636532395f244c5424696d706c2475323024247535622454247535642424475424313873706c69745f61745f756e636865636b65643137683765396534313435376636393734393145006e6578743c636f72653a3a736c6963653a3a697465723a3a497465723c636f72653a3a666d743a3a72743a3a506c616365686f6c6465723e3e007b696d706c2331377d005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542438697465725f6d75743137683030376635633136366631613761373245006172726179005f5a4e34636f7265337374723469746572323253706c6974496e7465726e616c244c5424502447542431346e6578745f696e636c75736976653137683938613230353930343932666138366445005f5a4e35325f244c542463686172247532302461732475323024636f72652e2e7374722e2e7061747465726e2e2e5061747465726e24475424313269735f7375666669785f6f663137683866653837336364343736333664316445005f5a4e34636f726533666d7439466f726d617474657238777261705f6275663137686636336162363038633262616362303045007b636c6f7375726523307d005f5a4e35365f244c54247573697a65247532302461732475323024636f72652e2e697465722e2e7472616974732e2e616363756d2e2e53756d244754243373756d3137683739356164323965353439386433333445005f5a4e34636f72653373747232315f244c5424696d706c2475323024737472244754243132636861725f696e64696365733137686466343535663065643137623532303045006765743c75382c207573697a653e005f5a4e34636f7265337074723132616c69676e5f6f66667365743137683534623332333739346162326331313545005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243961735f6368756e6b7331376831643562356538303063366463326238450061735f6368756e6b733c7573697a652c20343e005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243361646431376835666664656536393830656665666331450070616e69636b696e67006765745f756e636865636b65643c636f72653a3a666d743a3a72743a3a417267756d656e743e0064656275675f737472756374007b696d706c2332387d0065713c5b75385d2c205b75385d3e0044656275675475706c6500666d745f696e743c636f72653a3a666d743a3a6e756d3a3a55707065724865782c207536343e00636c616e67204c4c564d202872757374632076657273696f6e20312e37312e302d6e696768746c79202832663662633564323520323032332d30352d30392929006974657261746f72005f5a4e34636f726533737472313176616c69646174696f6e7331356e6578745f636f64655f706f696e74313768656364656330303032323838613566354500757466385f66697273745f627974650069735f636861725f626f756e64617279006d696e3c7573697a653e005f5a4e34636f72653373747235636f756e743330636f6e7461696e735f6e6f6e5f636f6e74696e756174696f6e5f627974653137686530636638653465356130663030393045005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137686134633765313364663063343439373145005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243361646431376833356564316564666234363437623138450077726974655f737472005f5a4e34636f726533666d74336e756d313247656e65726963526164697837666d745f696e743137686162643431393537653230363731373445006d617962655f756e696e697400696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e2c20636f72653a3a6f70733a3a72616e67653a3a52616e676546726f6d3c7573697a653e2c203132383e005f5a4e39395f244c5424636f72652e2e7374722e2e697465722e2e53706c6974496e636c7573697665244c54245024475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683536356238663563313134366339666645005f5a4e38315f244c5424636f72652e2e7374722e2e7061747465726e2e2e436861725365617263686572247532302461732475323024636f72652e2e7374722e2e7061747465726e2e2e53656172636865722447542431306e6578745f6d617463683137686231353436643361613035653433333145005f5a4e34636f72653463686172376d6574686f6473386c656e5f75746638313768343935363635353564666635366333654500656e636f64655f757466385f72617700616c6c6f6300747261697473005f5a4e34636f726535736c6963653469746572313349746572244c54245424475424336e65773137683436326338393130346236666239373745005f5a4e34636f7265336e756d32335f244c5424696d706c24753230247573697a652447542431327772617070696e675f6d756c3137683933396664623563663661656266303945006e6577006d656d6368720077726170005f5a4e34636f726533666d74336e756d313247656e65726963526164697837666d745f696e743137683330323730653937613764383866626145007061640070616e6963005f5a4e34636f726533666d74336e756d35335f244c5424696d706c2475323024636f72652e2e666d742e2e4c6f7765724865782475323024666f7224753230246936342447542433666d74313768663235653065383534373535336437314500696d7000616c7465726e617465006d6170005f5a4e3130325f244c5424636f72652e2e697465722e2e61646170746572732e2e6d61702e2e4d6170244c5424492443244624475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722447542434666f6c643137683439653563633739303661396231626645007772697465007b696d706c23377d006d696e5f62793c7573697a652c20666e28267573697a652c20267573697a6529202d3e20636f72653a3a636d703a3a4f72646572696e673e006765743c267374722c207573697a653e005f5a4e34636f726535736c69636535696e64657837345f244c5424696d706c2475323024636f72652e2e6f70732e2e696e6465782e2e496e646578244c542449244754242475323024666f72247532302424753562245424753564242447542435696e64657831376835623336343435386238326632343635450053706c6974496e7465726e616c006e6578743c636861723e0057726974650077726974655f636861723c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e007b696d706c2332367d005f5a4e34636f72653970616e69636b696e67313870616e69635f6e6f756e77696e645f666d743137683133386130386530383963323036303445005f5a4e34325f244c54242452462454247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d74313768633230363132656137383639386165344500666d74007b696d706c23307d004f7074696f6e007b696d706c23387d005f5a4e34636f726533707472376d75745f70747233315f244c5424696d706c2475323024244250246d757424753230245424475424336164643137686433383935323761353331303836366545006765745f756e636865636b65643c267374723e005f5a4e34636f726533666d7439466f726d6174746572313264656275675f73747275637431376838333134343030643138313466376534450070616e69635f737472005f5a4e34636f726533666d74386275696c64657273313564656275675f7475706c655f6e65773137683134383664383033383865636636373745005553495a455f4d41524b455200736c696365005f5a4e34636f7265336d656d377265706c6163653137683665313530623565366261663964346545007061645f696e74656772616c006765743c75383e005f5a4e34636f726535736c6963653469746572313349746572244c54245424475424336e65773137686231373834333338323430613463363745007b696d706c2331397d006e6578745f6d61746368005f5a4e34636f726536726573756c743139526573756c74244c542454244324452447542438616e645f7468656e3137686639613762303833656534636237383245005f5a4e37335f244c5424636f72652e2e666d742e2e6e756d2e2e5570706572486578247532302461732475323024636f72652e2e666d742e2e6e756d2e2e47656e657269635261646978244754243564696769743137683933663339316566393536306361643245005f5a4e34636f72653370747231303264726f705f696e5f706c616365244c542424524624636f72652e2e697465722e2e61646170746572732e2e636f706965642e2e436f70696564244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c542475382447542424475424244754243137683465633534623435323134663763393045005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683334323336653433336537396333623345006c74006368617273005f5a4e34636f72653373747232315f244c5424696d706c247532302473747224475424336765743137686361316261643162613538333362626645006765743c636f72653a3a6f70733a3a72616e67653a3a52616e6765546f3c7573697a653e3e00706f73745f696e635f73746172743c7573697a653e005f5a4e37355f244c54247573697a65247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c54242475356224542475356424244754242447542431336765745f756e636865636b65643137686630663432666234656339376261626145006164643c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e006d6574686f6473005f5a4e34636f726533666d74386275696c64657273313050616441646170746572347772617032385f24753762242475376224636c6f737572652475376424247537642431376862353032353031383864353564626337450063617061636974795f6f766572666c6f7700666d745f753634005f5a4e36385f244c5424636f72652e2e666d742e2e6275696c646572732e2e50616441646170746572247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f7374723137686539366438303337316562386433343445005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243361646431376836343831303738333031643161616237450049746572005f5a4e34636f72653373747232315f244c5424696d706c2475323024737472244754243563686172733137683635643537336338666664393434333645005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f723130616476616e63655f62793137683837343136383366376333383664636245006e6578745f636f64655f706f696e743c636f72653a3a736c6963653a3a697465723a3a497465723c75383e3e005f5a4e39335f244c5424636f72652e2e736c6963652e2e697465722e2e4368756e6b73244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137686264343939663734373230663065386245004f7264006164643c267374723e007b696d706c23367d005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f666d743137683565373464633863623261616161323645007b696d706c23327d005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542434697465723137686331616261316236653465646465623545005f5a4e34636f726533666d7439466f726d6174746572336e65773137686165623034366666366431666231663445005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243361646431376838353436653232346135313966363633450064656275675f7374727563745f6e657700746f5f7538005f5a4e34636f726533636d7035696d706c7336395f244c5424696d706c2475323024636f72652e2e636d702e2e5061727469616c4571244c54242452462442244754242475323024666f7224753230242452462441244754243265713137683436393566636435376362636161326145005f5a4e34636f726533666d743577726974653137683537653362636463656237646630393145006578706563745f6661696c6564006c656e5f6d69736d617463685f6661696c006f707300696e7472696e736963730073756d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e005f5a4e34636f7265336d656d377265706c61636531376838363534306363336630326138396663450069735f6e6f6e653c7573697a653e00697465723c5b7573697a653b20345d3e00696e746f5f697465723c5b7573697a653b20345d3e005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683366313636623661373436326234373945005f5a4e34636f726533666d7432727438417267756d656e7433666d74313768363232636537653835383430326338654500666d745f696e743c636f72653a3a666d743a3a6e756d3a3a4c6f7765724865782c207536343e00657175616c3c75382c2075383e005f5a4e34636f726535736c696365366d656d63687231326d656d6368725f6e616976653137686363623962373463393862393633336245006d656d6368725f6e6169766500616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23347d3a3a66696e6973683a3a7b636c6f737572655f656e7623307d3e005f5f616c6c6f635f6572726f725f68616e646c657200636f6e73745f707472005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f723373756d313768616537613566613764646461346162384500757466385f69735f636f6e745f62797465006e6578743c636f72653a3a666d743a3a72743a3a417267756d656e743e005f5a4e34636f726533666d74386275696c64657273313664656275675f7374727563745f6e65773137686135363836656238343531653037323245005f5a4e34636f72653970616e69636b696e67313370616e69635f646973706c6179313768663965353336303933393038663832624500656e64735f776974683c636861723e0065713c75382c2075383e007b696d706c23347d005f5a4e34636f726533737472313176616c69646174696f6e733137757466385f69735f636f6e745f6279746531376861396331376363326537313134623836450073706c69745f61745f756e636865636b65643c75383e0073706c69745f61743c75383e005f5a4e34636f72653373747235636f756e74313873756d5f62797465735f696e5f7573697a653137683733663965326535343130353136333245006e6578743c636f72653a3a666d743a3a72743a3a506c616365686f6c6465723e00417267756d656e74005f5a4e37355f244c54247573697a65247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c54242475356224542475356424244754242447542431336765745f756e636865636b6564313768656630633435353430343632353962624500636f6e7461696e735f7a65726f5f62797465005f5a4e37395f244c5424636f72652e2e726573756c742e2e526573756c74244c5424542443244524475424247532302461732475323024636f72652e2e6f70732e2e7472795f74726169742e2e54727924475424366272616e63683137683034646133323232663535363066313845005f5a4e34636f7265366f7074696f6e31336578706563745f6661696c65643137686332333330616533386638616564396545005f5a4e34636f726533707472376d75745f70747233315f244c5424696d706c2475323024244250246d7574247532302454244754243361646431376837336363316163653933303039363536450073756d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e2c207573697a653e005f5a4e35365f244c54247573697a65247532302461732475323024636f72652e2e697465722e2e7472616974732e2e616363756d2e2e53756d244754243373756d32385f24753762242475376224636c6f73757265247537642424753764243137683665653564323561643365666465373945007369676e5f61776172655f7a65726f5f70616400726561643c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e006e6578743c7573697a653e00756e777261705f6f723c267374723e005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243136616c69676e5f746f5f6f6666736574733137683265333033653231353164623038353745005f5a4e34636f726535736c69636532395f244c5424696d706c2475323024247535622454247535642424475424336765743137683037666466393631613031323632356145006e65773c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e007b696d706c2334347d0070616e69635f6e6f756e77696e645f666d740077726974655f7374723c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e577269746524475424313077726974655f636861723137683239666437616639333939643762333645005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243135636f70795f66726f6d5f736c69636531376c656e5f6d69736d617463685f6661696c3137686531663934356265353831313135613845006c6962726172792f616c6c6f632f7372632f6c69622e72732f402f616c6c6f632e643733613839653266303538366464312d6367752e30004974657261746f7200636f756e745f6368617273005f5a4e34636f72653469746572386164617074657273336d6170386d61705f666f6c6432385f24753762242475376224636c6f73757265247537642424753764243137686265643362346664336632356561633645005f5a4e34636f7265366f7074696f6e31354f7074696f6e244c542454244754243769735f6e6f6e653137683036303537623832613939663564313445005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542438616c69676e5f746f3137686361663565313535373365303734303345007b696d706c2331317d005f5a4e34636f726533636d70366d696e5f62793137683961363365346463336265666132393045005f5a4e34636f7265336d656d31326d617962655f756e696e697432304d61796265556e696e6974244c54245424475424357772697465313768643262633963366561386361383161624500656e636f64655f75746638005f5a4e34636f726533666d743557726974653977726974655f666d743137683364623431343565346436363932376245006669656c64005f5a4e36305f244c5424636f72652e2e63656c6c2e2e426f72726f774572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137686163386261333334363731373261333845006e6578743c75383e00746f5f7573697a65006d656d005f5a4e34636f7265337074723577726974653137683934303032343231393363646338316545005f5a4e38395f244c5424636f72652e2e6f70732e2e72616e67652e2e52616e6765244c54245424475424247532302461732475323024636f72652e2e697465722e2e72616e67652e2e52616e67654974657261746f72496d706c2447542439737065635f6e65787431376834303038636235396134653064623339450061735f7573697a65006164643c636f72653a3a666d743a3a72743a3a417267756d656e743e00696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e005f5a4e34636f7265336e756d32335f244c5424696d706c24753230247573697a652447542431327772617070696e675f73756231376838643635306338643866353735643162450069735f70726574747900616461707465727300726561643c636861723e007b696d706c23337d00636861725f696e646963657300616c69676e5f746f3c75382c207573697a653e007772617070696e675f6d756c0077726974653c75383e005f5a4e35305f244c5424753634247532302461732475323024636f72652e2e666d742e2e6e756d2e2e446973706c6179496e742447542435746f5f75383137683636316463333963356464386666653545007061747465726e0069735f7375666669785f6f66005f5a4e34636f726535736c696365366d656d63687231346d656d6368725f616c69676e6564313768643864383232303663636532343531614500526573756c740050616441646170746572005f5a4e34636f726533666d7439466f726d6174746572337061643137683433336537613934646232626438653245005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f7374723137683865303931326361326264646233386345005f5a4e34636f726533666d7432727431325553495a455f4d41524b455232385f24753762242475376224636c6f7375726524753764242475376424313768643137376134333532613130653633314500466e4f6e6365006e756d005f5a4e38315f244c5424636f72652e2e7374722e2e697465722e2e4368617273247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722447542435636f756e743137686638633866336432633063356164333545005f5a4e34636f726533666d7439466f726d617474657231397369676e5f61776172655f7a65726f5f7061643137683136323439616566366630343733333545006e65773c75383e007b696d706c23357d005f5a4e34636f726533636d70334f7264336d696e31376861623865636338303366663033636364450072756e005f5a4e34636f726533666d74386275696c64657273313044656275675475706c653969735f7072657474793137683131646663373739346165376162303045005f5a4e34636f726533666d7439466f726d617474657231327061645f696e74656772616c313277726974655f70726566697831376838346635386564303837613362643933450066756e6374696f6e00466f726d61747465720066696c746572006d61705f666f6c64005f5a4e38315f244c5424636f72652e2e7374722e2e697465722e2e4368617273247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683064323235303663643135633337363345007b696d706c2337307d005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683634663237353939353136663335636545005f5a4e35355f244c542424524624737472247532302461732475323024636f72652e2e7374722e2e7061747465726e2e2e5061747465726e24475424313269735f7375666669785f6f663137686536396533336230613062663235373545007772617070696e675f7375620077726974655f666d743c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e005f5a4e35616c6c6f63377261775f766563313763617061636974795f6f766572666c6f7731376837363964333737343539393364316265450063616c6c5f6f6e63653c636f72653a3a666d743a3a72743a3a5553495a455f4d41524b45523a3a7b636c6f737572655f656e7623307d2c2028267573697a652c20266d757420636f72653a3a666d743a3a466f726d6174746572293e0062000000020000000000740000003400000063617061636974795f6f766572666c6f77002f0000007261775f76656300590000005f5f72646c5f6f6f6d004f000000616c6c6f6300540000005f5f616c6c6f635f6572726f725f68616e646c65720000000000de1a0000020074000000cb2200006a01000077726974653c636861723e00c61e00006d617962655f756e696e6974007c2100006272616e63683c28292c20636f72653a3a666d743a3a4572726f723e00e90000006d75745f707472008a1f0000696e736572743c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e0003190000636f70795f6e6f6e6f7665726c617070696e673c75383e00b7040000466f726d617474657200752000007b696d706c2331377d00b01c0000737065635f6e6578743c7573697a653e0086190000706f73745f696e635f73746172743c7573697a653e00381800007b696d706c2332357d0057210000526573756c7400cb1d00006e6578745f636f64655f706f696e743c636f72653a3a736c6963653a3a697465723a3a497465723c75383e3e0034000000726561645f766f6c6174696c653c7573697a653e002b1a0000697465723c5b7573697a653b20345d3e00b91e00007265706c6163653c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e00711c00007b636c6f7375726523307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e00f719000073706c69745f61745f756e636865636b65643c75383e00ac1e00007265706c6163653c636861723e00701f000069735f6e6f6e653c7573697a653e00451a00006765743c267374722c207573697a653e00b02100007b696d706c2332367d00271e000069735f636861725f626f756e646172790038210000726573756c74008718000066756e6374696f6e00671c0000636f756e7400f00400007061645f696e74656772616c00111a0000616c69676e5f746f5f6f6666736574733c75382c207573697a653e008b1a00006c656e5f6d69736d617463685f6661696c00da0000006164643c75383e006e1900006e65773c75383e00e203000064696769740050180000666d743c28293e001f20000070616e69636b696e67007d1f0000756e777261705f6f723c267374723e00451d0000636f6e7461696e735f6e6f6e5f636f6e74696e756174696f6e5f6279746500cd000000616c69676e5f6f66667365743c75383e00bd1900006e65773c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e00d62000007b696d706c2331397d00102000007772617070696e675f73756200c9040000616c7465726e61746500fc1e00006c74003e1c00006d61705f666f6c6400511d000073756d5f62797465735f696e5f7573697a6500ae010000417267756d656e7400cb1e00004d61796265556e696e697400f4030000666d7400981f00006578706563745f6661696c6564009f1b0000636f6e7461696e735f7a65726f5f6279746500a911000072756e00a61d00007b696d706c2334347d006c1e00007b696d706c2332387d008d11000077726974655f707265666978008c180000466e4f6e636500d61a00006765743c267374723e005b000000636f6e73745f70747200971e00006e6578745f6d6174636800791a00006765743c75382c20636f72653a3a6f70733a3a72616e67653a3a52616e67653c7573697a653e3e00dd1e000077726974653c75383e00340100006164643c7573697a653e005d19000049746572003713000064656275675f7374727563745f6e6577004b1800007b696d706c2335337d00b30000006164643c636f72653a3a666d743a3a72743a3a417267756d656e743e00ed1c0000737472003d20000070616e69635f646973706c61793c267374723e00d0190000697465723c75383e00861a0000636f70795f66726f6d5f736c69636500271c00006d617000671e00007061747465726e00d9020000666d745f696e743c636f72653a3a666d743a3a6e756d3a3a4c6f7765724865782c207536343e00b015000066696e69736800dd0300007b696d706c2332397d0069210000616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23347d3a3a66696e6973683a3a7b636c6f737572655f656e7623307d3e003d210000756e777261705f6661696c656400201900006e6578743c75383e00931d000053706c6974496e7465726e616c00211d0000646f5f636f756e745f636861727300501900006e6578743c636f72653a3a666d743a3a72743a3a417267756d656e743e0011190000736c69636500c415000044656275675475706c65006c1c0000746f5f7573697a650062190000706f73745f696e635f73746172743c75383e005e1d000069746572000d1c000073756d00f71e00007b696d706c2335347d00931900007b696d706c2337307d00ca1a00006765745f756e636865636b65643c636f72653a3a666d743a3a72743a3a417267756d656e743e00841700007b696d706c23307d000f1d0000636861725f636f756e745f67656e6572616c5f6361736500841e000069735f7375666669785f6f6600311c0000666f6c643c7573697a652c20636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c207573697a652c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e007f100000777261705f6275663c636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23317d3a3a777261703a3a7b636c6f737572655f656e7623307d3e000918000077726974655f666d743c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e00e3010000666d745f753634002a000000636f7265001e1a000061735f6368756e6b733c7573697a652c20343e006211000064656275675f7475706c655f6669656c64315f66696e697368009c0100005553495a455f4d41524b455200221c0000616461707465727300f61f00007772617070696e675f6d756c00121c00007b636c6f7375726523307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e00331e00006765743c636f72653a3a6f70733a3a72616e67653a3a52616e6765546f3c7573697a653e3e00a60000006164643c5b7573697a653b20345d3e005b1c0000636f756e743c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e00ab190000696e746f5f697465723c5b7573697a653b20345d3e00c11b0000666f6c643c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a6d61703a3a6d61705f666f6c643a3a7b636c6f737572655f656e7623307d3c2675382c207573697a652c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e3e00e11600007b696d706c23317d005520000070616e69635f6e6f756e77696e645f666d7400902200006368617200511c000066696c74657200811c0000656e756d6572617465007b1b00006d656d6368725f6e6169766500e304000070616464696e6700160300007b696d706c2336347d00fc1b00007b696d706c2334387d00e61600007772617000f916000064656275675f7475706c655f6e657700431300007b696d706c23327d00b301000061735f7573697a6500011c000073756d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e00f21e0000696d706c7300f71b0000616363756d00071700005772697465002420000070616e696300441900006e6578743c636f72653a3a666d743a3a72743a3a506c616365686f6c6465723e000d1e0000636861727300821800006f707300952200006d6574686f6473005c1b000065713c75382c2075383e00ab1d00006e6578743c636861723e00ef0300007b696d706c2336357d00401e0000656e64735f776974683c636861723e00a71e00006d656d007f1e00007b696d706c23337d004920000070616e69635f73747200d61500006669656c6400381f00004f72640097010000727400de010000696d70008b1c00006e6578743c636f72653a3a736c6963653a3a697465723a3a497465723c636f72653a3a666d743a3a72743a3a506c616365686f6c6465723e3e00381900006e6578743c7573697a653e00b8190000497465724d757400c31100007772697465005f1a0000656e64735f776974683c75383e00c915000069735f707265747479002c1900006e6578743c5b7573697a653b20345d3e00e5020000666d745f696e743c636f72653a3a666d743a3a6e756d3a3a55707065724865782c207536343e00db1b0000616476616e63655f62793c636f72653a3a7374723a3a697465723a3a43686172496e64696365733e00d402000047656e657269635261646978004e1e0000747261697473008917000077726974655f7374723c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e00861d00006e65787400ce1b000073756d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e2c207573697a653e00981500007b696d706c23347d004813000077726974655f737472009a2200006c656e5f75746638001c1f000065713c5b75385d2c205b75385d3e005d010000726561643c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e00041a000073706c69745f61743c75383e00981d00006e6578745f696e636c75736976653c636861723e00040300007b696d706c2331317d0050010000726561643c636861723e00d907000070616400431c00007b636c6f7375726523307d3c2675382c207573697a652c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e00a217000077726974655f636861723c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e00d71d0000757466385f66697273745f6279746500391b00007b696d706c23357d00971c00006e6578743c636f72653a3a736c6963653a3a697465723a3a497465723c636f72653a3a666d743a3a72743a3a417267756d656e743e3e002b1f00006d696e5f62793c7573697a652c20666e28267573697a652c20267573697a6529202d3e20636f72653a3a636d703a3a4f72646572696e673e00591000006e657700df1f00006e756d007701000077726974653c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e00b41a0000696e646578005e1f00004f7074696f6e00631f000069735f736f6d653c7573697a653e00321300006275696c64657273001a1e0000636861725f696e6469636573007020000063656c6c00c00000006164643c267374723e00dd1900006765743c75382c207573697a653e00ef1a00007b696d706c23367d00251b00006765743c75383e00b51500007b636c6f7375726523307d00bf1d0000757466385f69735f636f6e745f6279746500bc1b00004974657261746f72009118000063616c6c5f6f6e63653c636f72653a3a666d743a3a72743a3a5553495a455f4d41524b45523a3a7b636c6f737572655f656e7623307d2c2028267573697a652c20266d757420636f72653a3a666d743a3a466f726d6174746572293e00871b00006d656d6368725f616c69676e656400ea190000616c69676e5f746f3c75382c207573697a653e00381a00006765745f756e636865636b65643c636f72653a3a666d743a3a72743a3a417267756d656e742c207573697a653e00410100006164643c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e00a61a0000697465725f6d75743c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e00591f00006f7074696f6e00a7220000656e636f64655f757466385f72617700ba1d000076616c69646174696f6e7300341b0000636d7000581e000067657400e21a00006765745f756e636865636b65643c267374723e00831100007b696d706c23377d001b1900007b696d706c233138317d00b71b00006974657261746f72007210000064656275675f73747275637400131b0000696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e2c20636f72653a3a6f70733a3a72616e67653a3a52616e676546726f6d3c7573697a653e3e00e81b00006e74683c636f72653a3a7374723a3a697465723a3a43686172496e64696365733e00b9220000656e636f64655f7574663800cf16000050616441646170746572006f1b00006d656d63687200531e00007b696d706c23387d00d7180000696e7472696e7369637300a2210000696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e2c20636f72653a3a6f70733a3a72616e67653a3a52616e676546726f6d3c7573697a653e2c203132383e00a61c000072616e676500902100007b696d706c2331357d00d60400007369676e5f61776172655f7a65726f5f70616400bc0400007369676e5f706c7573002f000000707472004100000064726f705f696e5f706c6163653c26636f72653a3a697465723a3a61646170746572733a3a636f706965643a3a436f706965643c636f72653a3a736c6963653a3a697465723a3a497465723c75383e3e3e00031d0000636f756e745f6368617273007a1900006e65773c5b7573697a653b20345d3e0070110000506f737450616464696e6700fb1d0000757466385f6163635f636f6e745f6279746500f41a0000696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e000a1f00007b696d706c23397d00b6110000676574636f756e74005c210000616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23347d3a3a6669656c643a3a7b636c6f737572655f656e7623307d3e004b1f00006d696e3c7573697a653e0009030000746f5f7538003e1b0000657175616c3c75382c2075383e008b210000617272617900000000000e00000002000000000074000000000000000e000000020074000000cb22000000000000412a000000726973637600012000000004100572763634693270305f6d3270305f613270305f633270300084000000040040000000010101fb0e0d0001010101000000010000016c6962726172792f616c6c6f632f73726300007261775f7665632e727300010000616c6c6f632e727300010000000009029a42010000000000038a040105050a030109020001090c000001010402000902a842010000000000038d0301050d0a030b09020001090c00000101ed1b0000040052030000010101fb0e0d0001010101000000010000016c6962726172792f636f72652f7372632f6f7073006c6962726172792f636f72652f7372632f707472006c6962726172792f636f72652f7372632f666d74006c6962726172792f636f72652f737263006c6962726172792f636f72652f7372632f736c6963652f69746572006c6962726172792f636f72652f7372632f697465722f747261697473006c6962726172792f636f72652f7372632f737472006c6962726172792f636f72652f7372632f69746572006c6962726172792f636f72652f7372632f697465722f6164617074657273006c6962726172792f636f72652f7372632f6d656d006c6962726172792f636f72652f7372632f6d6163726f73006c6962726172792f636f72652f7372632f736c696365006c6962726172792f636f72652f7372632f6e756d006c6962726172792f636f72652f7372632f6172726179006c6962726172792f636f72652f7372632f63686172000066756e6374696f6e2e7273000100006d6f642e72730002000072742e7273000300006e756d2e727300030000636f6e73745f7074722e727300020000696e7472696e736963732e7273000400006d75745f7074722e7273000200006d6f642e7273000300006d6163726f732e7273000500006974657261746f722e72730006000076616c69646174696f6e732e727300070000616363756d2e727300060000636d702e72730004000072616e67652e7273000800006d61702e72730009000066696c7465722e727300090000636f756e742e727300070000697465722e7273000700006d6f642e7273000a00006f7074696f6e2e7273000400006d6f642e7273000b00006d6f642e727300070000696e6465782e7273000c00007472616974732e7273000700006d6f642e7273000c000075696e745f6d6163726f732e7273000d0000697465722e7273000c000070616e69636b696e672e727300040000656e756d65726174652e72730009000063656c6c2e7273000400006275696c646572732e727300030000726573756c742e7273000400006d617962655f756e696e69742e7273000a00006d6f642e7273000e0000636d702e7273000c00007061747465726e2e7273000700006d656d6368722e7273000c00006d6574686f64732e7273000f000000000902747701000000000003f90101040205090a03860a090000010403050503d375090200010902000001010402000902787701000000000003ea030105010a03000900000109020000010104040009027a7701000000000003d2010105170a03130906000106039a7e0918000103e60109040001039a7e0924000105150603e80109020001051e0302090e00010405050d03b505091a00010406050903d20d090200010404051e03fa6c0904000104060509038613090400010405050d03ae72090800010406050903d20d090200010404051503fb6c09080001040605090385130902000106030009040001040405170603f56c0908000106039a7e0906000105140603f901090400010515030209040001051e037f091c000105150302090400010405050d03a305090200010406050903d20d090200010407050d039c73090c00010406050903e40c0902000106038f6b090a000104040514060381020902000105150301090400010407050d038b06090800010404051503f67909020001051e0302090a000105150301090200010405050d039905090400010406050903d20d090200010407050d039c73090c00010406050903e40c0902000106038f6b090800010407050d06038d08090400010404053e03827a09060001050d030209020001050a030109140001060b0300090200010904000001010408000902bc7801000000000003dd090105090a03e003091e0001051303a77c090c000106039b76090c000105090603f70d09040001051303ee7b0904000105190305090200010603967609020001050f0603fb0909020001050906030009020001038576090400010409051806038601090200010603fa7e09040001040a05150603b113090400010407050d03dc7409040001040b0505038c78090200010409051803ed0009080001040c051c03af7f090200010409051803d100090200010408050d03e50809020001050f031009020001050906030009020001052306030909020001051a06030009040001050906038d0409040001051a03f97b09020001051b03e90009020001053103a47f09060001051503dc000904000106038d7509060001050606039d0a09200001060b0300091c0001050003e3750904000104020509060394090926000106030009060001040805110603f900090400010402050903cd00090a000106030009040001040805110603b37f090400010603f3750914000105090603800b09020001040d05340353090600010408050d032e090400010603ff740910000105150603f30a090200010530030a0904000105230603000904000105300300090200010383750906000105090603800b090c0001040d0534035309040001040e050c039a7a090200010408050d039406090200010603ff74090c000105240603970a090a00010511030109040001030109140001050903fb7e090e0001040d053403bf01090800010408050d03c27e09080001051103fa00091000010603f175091000010603910a090200010301090400010603ee7509080001040d05340603d30a090200010906000001010408000902a07a01000000000003f2090105140a0301091c0001051103010904000105140302090e0001052c060300090200010b03000912000103897609040001050a0603f80909020001060b0300090a00010904000001010408000902f67a01000000000003bb0a01041405120a039b7a090200010408050c03e7050916000104150509039a78090200010408050c03e607090800010518030509040001051d060300090400010405050d0603dc7c09040001040a050903b87b09040001040b05000603a97d09120001041205260603910109040001051106030009020001040a05100603c70109040001040d053403fb0709040001040e050c039a7a090200010409051803997c09020001040b050d03a07f0904000105080301090800010516030a090400010505035b0904000105110306090400010508032109040001051a0305090400010505035a090400010511060300090200010505030009040001050c06032909040001051e030509040001051203010904000105050351090400010511060300090200010505030009040001050d06032f090400010412050903cb00090200010603f47e090400010409051806038601091e0001040b050d03a07f090400010508030109040001060359090400010603330908000106034d09040001050c06033b09040001050006034509040001051a060338090400010511035a0904000106030009040001051e06032e09040001051203010904000105050351090400010511060300090600010505030009040001050d06032f090200010412050903cb00090600010416050c03cc000904000105090304090200010417050c037d0904000104160513030f0904000104180509032c090800010603ec7d0904000104140603bc0709020001041803d87a090400010603ec7d0904000104140603bc07090200010603c4780902000104080603d40a0904000105120304090400010411050803c37509080001060365090400010409051806038601090200010603fa7e09040001040a05150603b113090400010407050d03dc7409040001040b0505038c78090200010409051803ed0009080001040c051c03af7f090200010409051803d100090200010402051f03bb0c0904000104190545036509060001051603800e090800010409051803e065090600010603fa7e09040001040a05150603b113090200010407050d03dc7409040001040b0505038c78090200010409051803ed0009080001040c051c03af7f090200010409051803d100090200010603fa7e090200010386010902000103fa7e09020001040a05150603b113090600010407050d03dc7409040001040b0505038c78090200010409051803ed0009080001040c051c03af7f090200010409051803d100090200010603fa7e09020001041105150603c7000922000105000603b97f09060001051b0603fe00090e00010534060300090400010533030009020001051b030009040001041a050d0603e7080902000104110505039a77090400010509035b09020001050c030609020001041b03e80a090200010603b874090200010419053806039908091200010405050d03867f090400010409051803e779090600010603fa7e09020001041105190603d0000904000105120301090200010507032309020001050606030009040001051203000902000106035d09020001050503230902000105110360090400010507032009020001050606030009040001051206035d090200010323090200010505060300090200010507030009040001050603000904000105120300090200010505030009020001051206035d0902000105050323090200010511036009020001050703200904000105060603000904000105120300090200010505030009020001040905180603120904000104110511034e09040001040905180332090200010603000906000103fa7e090400010386010904000103fa7e09040001038601090600010411051206035d090600010407050d03aa07090200010411050703e7780902000105060603000904000105120300090200010505030009020001040905180603120904000104110511035e09020001040905180322090200010603fa7e090400010411051b0603fe00090200010534060300090400010533030009020001051b030009040001041a050d0603e7080902000104110505039a7709040001050d0367090200010408051403f60909020001051b0317090400010535037009060001051503100904000106038d750906000103f30a09260001053006030a0904000105230603000904000105300300090200010383750906000105090603800b090e0001040d0534035309040001040e050c039a7a090200010408050d039406090200010603ff74090c000105280603e30a090a00010515030109040001050903b07e090e0001040d053403bf0109080001040e050c039a7a090400010408050d03a804090400010603eb7609100001040d05340603d30a0902000104080506031609040001060b030009140001090400000101041c0009026e7e01000000000003ed000105050a030709020001090c0000010104080009027c7e01000000000003b7080105090a03bb7909180001050b03c90609080001050903b77909040001050503c90609080001050e030e090200010409051803bc78090400010603fa7e0904000103860109040001040805150603cb0709220001051406030009020001051506030109020001052d0603000904000105150300090400010510060313090600010505060300090200010511060301090200010505060300090400010511060301090400010533036f09020001050503110904000105150304090200010505030f090600010403050c039978090600010603ed7e090a0001051d0603960109040001051b0603000902000103ea7e09020001040805090603eb080902000105190301090400010505030e090800010403050c039978090600010603ed7e090a0001051d0603960109040001051b0603000902000103ea7e09020001040805090603ec0809020001052d0307090400010405050d03ac7e090200010403050903eb7909040001051a060300090200010509030009020001040805110603cc07090400010409051803b078090200010408051d03b907091000010409051803c778090400010603fa7e0904000103860109080001040805150603bd0709120001051406030009020001051506030109020001052d060300090400010515030009040001040305090603c67809060001051a060300090200010509030009040001040805110603bc07090400010409051803c078090200010408051a03d707090a00010417050c03fc78090400010603a77e090600010408051a0603dd08090200010417050c03fc78090400010408051a038407090400010405050d03c27e090400010408050903bf0109040001052106030009040001050903000908000103a2770906000105020603e20809060001060b030009100001090400000101041e000902fa7f01000000000003ba0501040805090a03ba0609000001091200000101041e0009020c8001000000000003d50501040805090a039f060900000109120000010104200009021e8001000000000003f10c0105050a030109020001090c0000010104140009022c80010000000000038a0f01041c05050a038b7209020001090c00000101041c0009023a8001000000000003cf0001050e0a031009020001090c0000010104040009024880010000000000039901010407050d0a03f30609060001040405000603f3770908000106039301090800010421050903d602090200010404051403ea7c090400010603ad7f09080001052306032a0902000103e900090800010603ed7e090400010417050c0603ed03090a00010404050903817d090a0001050e032e09160001060b0300090200010417050d0603d20209040001090e00000101041f000902b880010000000000031e010412050c0a03ce040946000104190523039c0d091800010423050d03d26e09040001041f034a090a00010301090400010412050c03c704090e00010424051903b17e090800010417050c0342090a00010425050803cb7d09080001050b030d0906000106034809040001050c0603390902000105090304090c0001050b037b090200010402051f03890d09060001051b03010908000104250508039273090400010603ac7f090e000105100603eb00090600010405050d03b406090400010425051503c679090400010529030409060001041a050d03e508090200010425050503c67609020001051503d2000908000105290304090a0001041a050d03e408090200010425050503c67609020001050903db0009080001050b037209020001050c03580906000105090304090c0001050b037b09020001060348090400010603e1000904000106039f7f09040001050c06033909060001050b037f090c000106034809080001042405200603b403090200010511060300090200010417050c0603ac7f090800010423050d03fb7d090200010424051c03dd02090400010603c87c09040001041f051006032109140001051103010906000106035e090e00010419050906038912090800010603f76d09040001041f050606032a09100001060b0300091a00010904000001010408000902748201000000000003a20101052b0a0301090c00010426050803f60b09020001050d031f09040001050f0363090800010513032009060001050d06030009040001051206030109080001050d06030009040001050f060361090c00010513032209060001050d06030009040001051206030109080001050d06030009060001051206030109080001050d060300090400010512060303090c0001050d06030009060001051206030109080001050d06030009060001051206030109080001050d06030009060001051206030109080001050d06030009040001040805090603dc73090a000105060301090a0001060b0300090200010904000001010408000902288301000000000003be010105090a0301090200010506030109300001060b0300090200010904000001010408000902608301000000000003c5010105090a030109000001090a0000010104080009026a8301000000000003c9010105090a030109020001052b0359090c00010426050803f60b09020001050d031f09040001050f0363090800010513032009060001050d06030009040001051206030109080001050d06030009040001050f060361090c00010513032209060001050d06030009040001051206030109080001050d06030009060001051206030109080001050d060300090400010512060303090c0001050d06030009060001051206030109080001050d06030009060001051206030109080001050d06030009060001051206030109080001050d06030009040001040805090603dc73090a000105060328090a0001060b0300090200010904000001010408000902208401000000000003cd010105090a0301090200010371091e00010506031009140001060b030009020001090400000101041f0009025a8401000000000003b3020105170a0301091200010420050903f10709040001041f03a078090200010603ba7d0908000105100603b602090400010408050903c10b09040001041f050006038972090400010408050903f70d09040001041f05100603bf740904000105000603ca7d09020001051e0603c002090400010603c07d0904000105140603b702090a00010408050903be0909040001041f051503c376091600010603c87d09020001040805090603f50b090e0001041f051e03cb76090a00010408050903b50909020001042003a70309040001041f051103a673090200010408051403e406090c00010603da7609040001041f05210603bb02090200010408051703e806090400010414050903f002090800010408051303947d090a0001051403010904000103010904000105180301090800010509037709080001041f0511039c79091400010408050903e40609040001041f0511039c79090a00010408050903b80909080001041f050006038b740912000105090603b502090200010311090400010506030209060001060b03000910000109040000010104080009027a8501000000000003e40f0105090a03907c090c0001041f050503a376090c00010408050903cf0d090c0001041f050c03fd72090e0001050006039c7d09020001050c03e40209040001039c7d09020001042005090603a60a09020001041f051403c07809020001050006039a7d090a0001051403e60209020001040805090603910b09080001041f051403ef740906000104080509038f0909020001041f051503f2760914000104080509038e0909020001041f03f776091600010408050603fd0c09040001060b0300090a000109040000010104190009021286010000000000038a1a01050d0a030109020001090c000001010408000902208601000000000003cf110105090a03ec01090000010916000001010422000902368601000000000003820101040805090a03f20a090a00010422051e038f75090200010408050903f10a09020001041f050503a376091000010408050903cf0d090c0001041f050c03fd7209140001050006039c7d09020001050c03e40209040001039c7d09020001042005090603a60a09020001041f051403c07809020001050006039a7d090a0001051403e60209020001040805090603910b09080001041f051403ef740906000104080509038f0909020001041f051503f2760914000104080509038e0909020001041f03f776091600010422050f03977e09040001060b0300090800010904000001010404000902d886010000000000039901010407050d0a03f30609060001040405000603f3770908000106039401090800010421050903d502090200010404051403ea7c090400010603ad7f09080001052306032a0902000103ea00090800010603ec7e090400010417050c0603ed03090a00010404050903817d090a0001050e032e09160001060b0300090200010417050d0603d20209040001090e00000101004743433a2028292031322e322e30004c696e6b65723a204c4c442031362e302e320000000000000000000000000000000000000000000000000000000000010000000400f1ff000000000000000000000000000000000000000000000300ea2601000000000000000000000000000000000000000300ee2601000000000000000000000000000000000000000300222701000000000000000000000000001e00000000000300222701000000000000000000000000002a0000000100050008bd01000000000010000000000000005300000002000300aa880100000000004e000000000000009b0000000000030020280100000000000000000000000000a70000000100010091040100000000000c00000000000000d30000000000030064280100000000000000000000000000df000000000003008e280100000000000000000000000000eb00000002000300ca7401000000000036000000000000004501000002000300ae91010000000000080000000000000054010000020003000c950100000000002800000000000000cd010000000003007e290100000000000000000000000000d901000000000300ac290100000000000000000000000000e501000000000300d4290100000000000000000000000000f1010000020003009c7201000000000022000000000000006c02000002000300c86f010000000000d6000000000000000003000002000300be720100000000003a000000000000003903000002000300f47301000000000042000000000000007803000000000300722a010000000000000000000000000084030000000003009c2a01000000000000000000000000009003000002000300f872010000000000fc0000000000000018040000020003003a7201000000000062000000000000004b04000000000300e82b0100000000000000000000000000570400000100010056040100000000000c000000000000008204000000000300082c01000000000000000000000000008f040000010001004c040100000000000a00000000000000ba04000002000300ce710100000000006c00000000000000ed04000002000300dc90010000000000ba000000000000006e05000002000300fa8c0100000000005400000000000000af05000002000300c08f010000000000a2000000000000004c06000002000300308a0100000000005600000000000000ab060000000003009a2e0100000000000000000000000000b8060000010001009d040100000000001100000000000000e406000000000300de2e0100000000000000000000000000f106000000000300082f0100000000000000000000000000fe06000000000300982f01000000000000000000000000000b07000000000300c62f01000000000000000000000000001807000000000300ee2f010000000000000000000000000025070000000003008c3001000000000000000000000000003207000000000300b63001000000000000000000000000003f0700000200030012860100000000000e00000000000000a50700000000030064320100000000000000000000000000b20700000100010070040100000000002100000000000000bb070000020003006e7e0100000000000e00000000000000e807000002000300d09101000000000072000000000000006908000002000300fc750100000000006001000000000000a5080000020003004e8d0100000000007c01000000000000eb0800000200030098960100000000008605000000000000200900000200030000750100000000007a000000000000006109000002000300be430100000000005800000000000000b8090000020003000e430100000000005800000000000000140a000002000300664301000000000058000000000000006e0a00000200030068a30100000000008601000000000000af0a00000200030034950100000000006401000000000000e90a00000200030012450100000000005800000000000000480b000002000300b6420100000000005800000000000000a30b000002000300369f0100000000009200000000000000de0b000000000300943b0100000000000000000000000000eb0b00000100010040090100000000001c00000000000000f50b0000000003002e3c0100000000000000000000000000020c00000100010060090100000000002b000000000000002d0c000000000300363c01000000000000000000000000003a0c00000100010018020100000000002000000000000000650c000000000300403c0100000000000000000000000000720c000000000300483c01000000000000000000000000007f0c0000020003001e800100000000000e00000000000000b20c000002000300c89f010000000000a003000000000000f60c000002000300164401000000000052000000000000004f0d0000020003006a450100000000004e00000000000000a20d00000200030068440100000000005800000000000000f50d000002000300c0440100000000005200000000000000550e0000020003001e9c01000000000018030000000000008c0e00000000030014400100000000000000000000000000990e0000000003001c400100000000000000000000000000a60e000001000100b0090100000000002000000000000000d10e00000000030062410100000000000000000000000000de0e0000000003006a410100000000000000000000000000eb0e000001000100b0010100000000002000000000000000150f00000000030074410100000000000000000000000000220f0000000003007c4101000000000000000000000000002f0f0000000003008e4101000000000000000000000000003c0f00000000030096410100000000000000000000000000490f000000000300a0410100000000000000000000000000560f000000000300a8410100000000000000000000000000630f000000000300b2410100000000000000000000000000700f00000100010050070100000000002b000000000000009a0f000000000300c2410100000000000000000000000000a70f000001000100d0010100000000001c00000000000000ad0f000000000300cc410100000000000000000000000000ba0f000001000100f0010100000000002100000000000000c00f000000000300d8410100000000000000000000000000cd0f000000000300e4410100000000000000000000000000da0f000000000300f0410100000000000000000000000000000000000000030002420100000000000000000000000000e70f00000200030002420100000000000a00000000000000000000000000030002420100000000000000000000000000f90f0000020003005c77010000000000180000000000000000000000000003000c4201000000000000000000000000002e100000020003000c42010000000000080000000000000000000000000003000c42010000000000000000000000000039100000020003000268010000000000d403000000000000000000000000030014420100000000000000000000000000c41000000200030014420100000000000800000000000000000000000000030014420100000000000000000000000000d110000002000300d66b010000000000f20300000000000000000000000003001c4201000000000000000000000000005e110000020003001c420100000000004e0000000000000000000000000003001c42010000000000000000000000000000000000000003001e42010000000000000000000000000000000000000003002842010000000000000000000000000000000000000003006a4201000000000000000000000000006b110000020003006a42010000000000300000000000000000000000000003006a42010000000000000000000000000000000000000003006c42010000000000000000000000000000000000000003007242010000000000000000000000000000000000000003009a4201000000000000000000000000007d110000020003009a420100000000000e0000000000000000000000000003009a42010000000000000000000000000000000000000003009a42010000000000000000000000000000000000000003009a42010000000000000000000000000000000000000003009c42010000000000000000000000000000000000000003009c42010000000000000000000000000000000000000003009e420100000000000000000000000000b6110000020003003a800100000000000e000000000000000000000000000300a84201000000000000000000000000000000000000000300a8420100000000000000000000000000f111000002000300a8420100000000000e000000000000000000000000000300a84201000000000000000000000000000000000000000300a84201000000000000000000000000000000000000000300a84201000000000000000000000000000000000000000300aa4201000000000000000000000000000000000000000300aa4201000000000000000000000000000000000000000300ac4201000000000000000000000000000000000000000300b64201000000000000000000000000000000000000000300b64201000000000000000000000000000000000000000300b64201000000000000000000000000000000000000000300b84201000000000000000000000000000000000000000300bc420100000000000000000000000000fb11000000000300ee4201000000000000000000000000000812000000000300f642010000000000000000000000000000000000000003000e43010000000000000000000000000000000000000003000e43010000000000000000000000000000000000000003001043010000000000000000000000000000000000000003001443010000000000000000000000000015120000000003004643010000000000000000000000000022120000000003004e43010000000000000000000000000000000000000003006643010000000000000000000000000000000000000003006643010000000000000000000000000000000000000003006843010000000000000000000000000000000000000003006c4301000000000000000000000000002f120000000003009e4301000000000000000000000000003c12000000000300a64301000000000000000000000000000000000000000300be4301000000000000000000000000000000000000000300be4301000000000000000000000000000000000000000300c04301000000000000000000000000000000000000000300c44301000000000000000000000000004912000000000300f64301000000000000000000000000005612000000000300fe43010000000000000000000000000000000000000003001644010000000000000000000000000000000000000003001644010000000000000000000000000000000000000003001844010000000000000000000000000000000000000003001a4401000000000000000000000000006312000002000300428f0100000000007e00000000000000e81200000000030048440100000000000000000000000000f5120000000003005044010000000000000000000000000000000000000003006844010000000000000000000000000000000000000003006844010000000000000000000000000000000000000003006a44010000000000000000000000000000000000000003006e4401000000000000000000000000000213000000000300a04401000000000000000000000000000f13000000000300a84401000000000000000000000000000000000000000300c04401000000000000000000000000000000000000000300c04401000000000000000000000000000000000000000300c24401000000000000000000000000000000000000000300c44401000000000000000000000000001c13000002000300ca8e0100000000007800000000000000a213000000000300f2440100000000000000000000000000af13000000000300fa440100000000000000000000000000000000000000030012450100000000000000000000000000000000000000030012450100000000000000000000000000000000000000030014450100000000000000000000000000000000000000030018450100000000000000000000000000bc130000000003004a450100000000000000000000000000c9130000000003005245010000000000000000000000000000000000000003006a45010000000000000000000000000000000000000003006a45010000000000000000000000000000000000000003006c450100000000000000000000000000000000000000030070450100000000000000000000000000d61300000000030096450100000000000000000000000000e3130000000003009e4501000000000000000000000000000000000000000300b8450100000000000000000000000000f013000002000300b8450100000000009a000000000000000000000000000300b84501000000000000000000000000000000000000000300ba4501000000000000000000000000000000000000000300c24501000000000000000000000000003614000000000300d845010000000000000000000000000043140000010001003802010000000000400000000000000000000000000003005246010000000000000000000000000081140000020003005246010000000000dc00000000000000000000000000030052460100000000000000000000000000000000000000030056460100000000000000000000000000000000000000030062460100000000000000000000000000c3140000020003002e47010000000000ee1a00000000000000000000000003002e4701000000000000000000000000000715000000000400f0bb01000000000000000000000000001115000000000400f8bb01000000000000000000000000001b1500000000040000bc0100000000000000000000000000251500000000040008bc01000000000000000000000000002f1500000000040010bc0100000000000000000000000000391500000000040018bc0100000000000000000000000000431500000000040020bc01000000000000000000000000004d1500000000040028bc010000000000000000000000000000000000000003002e47010000000000000000000000000000000000000003003047010000000000000000000000000000000000000003004a4701000000000000000000000000005715000000000300ca4701000000000000000000000000006415000000000300de47010000000000000000000000000071150000000003002a4801000000000000000000000000007e150000000003003e4801000000000000000000000000008b15000000000300884801000000000000000000000000009815000000000300a2480100000000000000000000000000a515000000000300e8480100000000000000000000000000b215000000000300fe48010000000000000000000000000000000000000003001c620100000000000000000000000000bf150000020003001c62010000000000140400000000000000000000000003001c62010000000000000000000000000000000000000003001e620100000000000000000000000000000000000000030038620100000000000000000000000000011600000200030030660100000000003c000000000000003b16000000000300fe620100000000000000000000000000481600000100010060030100000000001c00000000000000511600000200030076660100000000004c000000000000008a16000002000300c2660100000000004c00000000000000d5160000020003002c800100000000000e0000000000000008170000000003007665010000000000000000000000000015170000000003008a6501000000000000000000000000002217000000000300946501000000000000000000000000002f170000000003009e6501000000000000000000000000003c17000000000300a86501000000000000000000000000004917000001000100000301000000000021000000000000005217000000000300b26501000000000000000000000000005f17000001000100300301000000000024000000000000006817000000000300c06501000000000000000000000000007517000000000300ca6501000000000000000000000000008217000001000100d00201000000000021000000000000008b17000000000300d46501000000000000000000000000009817000000000300de650100000000000000000000000000a517000000000300e8650100000000000000000000000000b217000001000100a0020100000000002300000000000000bb17000000000300f6650100000000000000000000000000c817000001000100a0030100000000001000000000000000f317000000000300106601000000000000000000000000000018000001000100e80301000000000010000000000000002b180000020003006c660100000000000a000000000000006118000000000300226601000000000000000000000000000000000000000300306601000000000000000000000000000000000000000300306601000000000000000000000000006e18000000000300486601000000000000000000000000007b180000000003005666010000000000000000000000000000000000000003006c66010000000000000000000000000000000000000003006c66010000000000000000000000000000000000000003007666010000000000000000000000000000000000000003007666010000000000000000000000000088180000000003009466010000000000000000000000000095180000000003009e660100000000000000000000000000a218000000000300ac6601000000000000000000000000000000000000000300c26601000000000000000000000000000000000000000300c2660100000000000000000000000000af18000000000300e2660100000000000000000000000000bc18000000000300ec660100000000000000000000000000c91800000000030002670100000000000000000000000000d618000001000100f8030100000000000d0000000000000000000000000003000e67010000000000000000000000000001190000020003000e67010000000000f40000000000000000000000000003000e6701000000000000000000000000004019000000000300da6701000000000000000000000000004d19000000000300ee6701000000000000000000000000005a19000000000300f867010000000000000000000000000000000000000003000268010000000000000000000000000000000000000003000268010000000000000000000000000000000000000003000468010000000000000000000000000000000000000003001c680100000000000000000000000000671900000000030022680100000000000000000000000000741900000100050060bc010000000000a80000000000000098190000000003002e680100000000000000000000000000a519000000000300d8690100000000000000000000000000b3190000000003001a6a0100000000000000000000000000c1190000000003004a6b0100000000000000000000000000cf19000000000300546b0100000000000000000000000000dd19000000000300626b0100000000000000000000000000eb19000000000300766b0100000000000000000000000000f919000000000300806b0100000000000000000000000000061a000000000300946b0100000000000000000000000000131a0000000003009c6b0100000000000000000000000000211a000001000100780201000000000020000000000000004b1a000000000300a66b0100000000000000000000000000581a000000000300ae6b0100000000000000000000000000651a000000000300b86b0100000000000000000000000000731a000000000300c06b01000000000000000000000000000000000000000300d66b01000000000000000000000000000000000000000300d66b01000000000000000000000000000000000000000300d86b01000000000000000000000000000000000000000300f26b0100000000000000000000000000811a000000000300f26b01000000000000000000000000008f1a000000000300106c01000000000000000000000000009d1a0000000003005c6c0100000000000000000000000000ab1a000000000300046d0100000000000000000000000000b91a000000000300546f0100000000000000000000000000c71a0000000003005e6f0100000000000000000000000000d51a0000000003006c6f0100000000000000000000000000e31a000000000300806f0100000000000000000000000000f11a000000000300986f0100000000000000000000000000ff1a000000000300a06f01000000000000000000000000000d1b000000000300aa6f01000000000000000000000000001b1b000000000300b26f01000000000000000000000000000000000000000300c86f01000000000000000000000000000000000000000300c86f01000000000000000000000000000000000000000300ca6f01000000000000000000000000000000000000000300d86f0100000000000000000000000000291b0000020003009e700100000000005200000000000000711b000002000300f0700100000000003400000000000000cb1b0000000003007c700100000000000000000000000000d91b0000010001001004010000000000190000000000000000000000000003009e70010000000000000000000000000000000000000003009e7001000000000000000000000000000000000000000300a07001000000000000000000000000000000000000000300a6700100000000000000000000000000e21b000002000300a6910100000000000800000000000000ef1b000002000300c6910100000000000a000000000000000000000000000300f07001000000000000000000000000000000000000000300f07001000000000000000000000000000000000000000300f27001000000000000000000000000000000000000000300f47001000000000000000000000000000a1c0000020003002471010000000000740000000000000000000000000003002471010000000000000000000000000000000000000003002471010000000000000000000000000000000000000003002671010000000000000000000000000000000000000003002c710100000000000000000000000000551c00000200030018880100000000006200000000000000000000000000030098710100000000000000000000000000881c0000020003009871010000000000360000000000000000000000000003009871010000000000000000000000000000000000000003009a71010000000000000000000000000000000000000003009c7101000000000000000000000000000000000000000300ce7101000000000000000000000000000000000000000300ce7101000000000000000000000000000000000000000300d07101000000000000000000000000000000000000000300dc71010000000000000000000000000000000000000003003a72010000000000000000000000000000000000000003003a72010000000000000000000000000000000000000003003c72010000000000000000000000000000000000000003004872010000000000000000000000000000000000000003009c72010000000000000000000000000000000000000003009c7201000000000000000000000000000000000000000300be7201000000000000000000000000000000000000000300be7201000000000000000000000000000000000000000300c07201000000000000000000000000000000000000000300c67201000000000000000000000000000000000000000300f87201000000000000000000000000000000000000000300f87201000000000000000000000000000000000000000300fa720100000000000000000000000000000000000000030008730100000000000000000000000000d51c00000000030024730100000000000000000000000000e31c00000100010062040100000000000b000000000000000f1d000000000300807301000000000000000000000000001d1d000000000300da7301000000000000000000000000000000000000000300f47301000000000000000000000000000000000000000300f47301000000000000000000000000000000000000000300367401000000000000000000000000002b1d0000020003003674010000000000920000000000000000000000000003003674010000000000000000000000000000000000000003003874010000000000000000000000000000000000000003003a740100000000000000000000000000861d0000000003003e740100000000000000000000000000941d000000000100600101000000000000000000000000009e1d0000000003004c740100000000000000000000000000a71d00000000030052740100000000000000000000000000b51d0000010001002b050100000000000f00000000000000e01d0000000003005e740100000000000000000000000000e91d00000000030064740100000000000000000000000000f71d00000100010020050100000000000b00000000000000221e000000000300707401000000000000000000000000002b1e00000000030074740100000000000000000000000000391e000001000100f0040100000000000f00000000000000641e0000000003007c740100000000000000000000000000721e000001000100000501000000000020000000000000009d1e00000000030088740100000000000000000000000000a61e0000000003008e740100000000000000000000000000b41e0000000003009e740100000000000000000000000000bd1e000000000300a2740100000000000000000000000000cb1e000001000100ae040100000000000700000000000000f61e000000000300aa740100000000000000000000000000041f000001000100b80401000000000020000000000000002f1f0000020003007a8501000000000098000000000000000000000000000300c8740100000000000000000000000000751f000002000300c87401000000000002000000000000000000000000000300c87401000000000000000000000000000000000000000300ca7401000000000000000000000000000000000000000300ca74010000000000000000000000000000000000000003000075010000000000000000000000000000000000000003000075010000000000000000000000000000000000000003000275010000000000000000000000000000000000000003000675010000000000000000000000000000000000000003007a750100000000000000000000000000b41f0000020003007a75010000000000820000000000000000000000000003007a75010000000000000000000000000000000000000003007c7501000000000000000000000000000000000000000300807501000000000000000000000000000000000000000300fc7501000000000000000000000000000000000000000300fc75010000000000000000000000000000000000000003000076010000000000000000000000000000000000000003002476010000000000000000000000000000000000000003005c77010000000000000000000000000000000000000003005c770100000000000000000000000000000000000000030074770100000000000000000000000000f51f0000020003007477010000000000040000000000000000000000000003007477010000000000000000000000000000000000000003007477010000000000000000000000000000000000000003007477010000000000000000000000000000000000000003007477010000000000000000000000000000000000000003007677010000000000000000000000000000000000000003007677010000000000000000000000000000000000000003007877010000000000000000000000000000000000000003007877010000000000000000000000000000000000000003007877010000000000000000000000000030200000020003007877010000000000020000000000000000000000000003007877010000000000000000000000000000000000000003007877010000000000000000000000000000000000000003007877010000000000000000000000000000000000000003007877010000000000000000000000000000000000000003007a77010000000000000000000000000000000000000003007a770100000000000000000000000000ba2000000000040030bc0100000000000000000000000000c4200000020003007a77010000000000420100000000000000000000000003007a77010000000000000000000000000000000000000003007a77010000000000000000000000000000000000000003007a77010000000000000000000000000000000000000003007c77010000000000000000000000000000000000000003007e770100000000000000000000000000000000000000030080770100000000000000000000000000f5200000000003008c77010000000000000000000000000003210000010001009e05010000000000c80000000000000000000000000003009877010000000000000000000000000000000000000003009c7701000000000000000000000000002f21000000000300a07701000000000000000000000000000000000000000300c07701000000000000000000000000000000000000000300c27701000000000000000000000000000000000000000300d07701000000000000000000000000000000000000000300ea7701000000000000000000000000000000000000000300ea7701000000000000000000000000000000000000000300ec7701000000000000000000000000000000000000000300ec7701000000000000000000000000000000000000000300f07701000000000000000000000000000000000000000300f07701000000000000000000000000000000000000000300f47701000000000000000000000000000000000000000300f47701000000000000000000000000000000000000000300fc7701000000000000000000000000000000000000000300fc7701000000000000000000000000000000000000000300fe7701000000000000000000000000000000000000000300fe77010000000000000000000000000000000000000003000678010000000000000000000000000000000000000003000678010000000000000000000000000000000000000003000878010000000000000000000000000000000000000003000878010000000000000000000000000000000000000003000c78010000000000000000000000000000000000000003000c78010000000000000000000000000000000000000003001478010000000000000000000000000000000000000003001478010000000000000000000000000000000000000003001a78010000000000000000000000000000000000000003001e78010000000000000000000000000000000000000003002278010000000000000000000000000000000000000003003e78010000000000000000000000000000000000000003004278010000000000000000000000000000000000000003004478010000000000000000000000000000000000000003004478010000000000000000000000000000000000000003004678010000000000000000000000000000000000000003004678010000000000000000000000000000000000000003005278010000000000000000000000000000000000000003005278010000000000000000000000000000000000000003005478010000000000000000000000000000000000000003005478010000000000000000000000000000000000000003005e78010000000000000000000000000000000000000003005e78010000000000000000000000000000000000000003006078010000000000000000000000000000000000000003006478010000000000000000000000000000000000000003006c78010000000000000000000000000000000000000003006c78010000000000000000000000000000000000000003006e78010000000000000000000000000000000000000003006e78010000000000000000000000000000000000000003007878010000000000000000000000000000000000000003007a78010000000000000000000000000000000000000003007e78010000000000000000000000000000000000000003007e78010000000000000000000000000000000000000003008078010000000000000000000000000000000000000003008078010000000000000000000000000000000000000003008c78010000000000000000000000000000000000000003008c78010000000000000000000000000000000000000003008e78010000000000000000000000000000000000000003008e78010000000000000000000000000000000000000003009678010000000000000000000000000000000000000003009678010000000000000000000000000000000000000003009a78010000000000000000000000000000000000000003009a7801000000000000000000000000000000000000000300a07801000000000000000000000000000000000000000300a07801000000000000000000000000003d21000000000300a27801000000000000000000000000004b21000001000100600901000000000000000000000000000000000000000300a27801000000000000000000000000007621000002000300bc78010000000000e4010000000000000000000000000300b67801000000000000000000000000000000000000000300b87801000000000000000000000000000000000000000300bc7801000000000000000000000000000000000000000300bc7801000000000000000000000000000000000000000300bc7801000000000000000000000000000000000000000300bc7801000000000000000000000000000000000000000300bc7801000000000000000000000000000000000000000300be7801000000000000000000000000000000000000000300d87801000000000000000000000000000000000000000300da7801000000000000000000000000000000000000000300da7801000000000000000000000000000000000000000300e67801000000000000000000000000000000000000000300e67801000000000000000000000000000000000000000300f27801000000000000000000000000000000000000000300f67801000000000000000000000000000000000000000300f67801000000000000000000000000000000000000000300fa7801000000000000000000000000000000000000000300fa7801000000000000000000000000000000000000000300fc7801000000000000000000000000000000000000000300fe78010000000000000000000000000000000000000003000079010000000000000000000000000000000000000003000279010000000000000000000000000000000000000003000679010000000000000000000000000000000000000003000879010000000000000000000000000000000000000003000879010000000000000000000000000000000000000003000c79010000000000000000000000000000000000000003000c79010000000000000000000000000000000000000003001079010000000000000000000000000000000000000003001479010000000000000000000000000000000000000003001479010000000000000000000000000000000000000003001679010000000000000000000000000000000000000003001679010000000000000000000000000000000000000003001e79010000000000000000000000000000000000000003001e79010000000000000000000000000000000000000003002079010000000000000000000000000000000000000003002079010000000000000000000000000000000000000003002279010000000000000000000000000000000000000003002279010000000000000000000000000000000000000003002479010000000000000000000000000000000000000003002479010000000000000000000000000000000000000003002679010000000000000000000000000000000000000003002879010000000000000000000000000000000000000003002a79010000000000000000000000000000000000000003002e79010000000000000000000000000000000000000003003279010000000000000000000000000000000000000003003279010000000000000000000000000000000000000003003479010000000000000000000000000000000000000003003479010000000000000000000000000000000000000003003679010000000000000000000000000000000000000003003679010000000000000000000000000000000000000003003c79010000000000000000000000000000000000000003003c790100000000000000000000000000000000000000030040790100000000000000000000000000000000000000030040790100000000000000000000000000000000000000030046790100000000000000000000000000000000000000030046790100000000000000000000000000af21000002000300a07a01000000000056000000000000000000000000000300667901000000000000000000000000000000000000000300827901000000000000000000000000000000000000000300867901000000000000000000000000000000000000000300ac7901000000000000000000000000000000000000000300ac7901000000000000000000000000000000000000000300b27901000000000000000000000000000000000000000300b27901000000000000000000000000000000000000000300b67901000000000000000000000000000000000000000300b67901000000000000000000000000000000000000000300c07901000000000000000000000000000000000000000300c07901000000000000000000000000000000000000000300c47901000000000000000000000000000000000000000300c47901000000000000000000000000000000000000000300c87901000000000000000000000000000000000000000300c87901000000000000000000000000000000000000000300dc7901000000000000000000000000000000000000000300de7901000000000000000000000000000000000000000300de7901000000000000000000000000000000000000000300e47901000000000000000000000000000000000000000300e47901000000000000000000000000000000000000000300e87901000000000000000000000000000000000000000300e87901000000000000000000000000000000000000000300f87901000000000000000000000000000000000000000300f87901000000000000000000000000000000000000000300fa7901000000000000000000000000000000000000000300fa7901000000000000000000000000000000000000000300fe7901000000000000000000000000000000000000000300027a01000000000000000000000000000000000000000300047a010000000000000000000000000000000000000003000a7a01000000000000000000000000000000000000000300167a010000000000000000000000000000000000000003001a7a010000000000000000000000000000000000000003001a7a010000000000000000000000000000000000000003001c7a010000000000000000000000000000000000000003001c7a010000000000000000000000000000000000000003001e7a010000000000000000000000000000000000000003001e7a010000000000000000000000000000000000000003002a7a010000000000000000000000000000000000000003002a7a01000000000000000000000000000000000000000300347a01000000000000000000000000000000000000000300387a010000000000000000000000000000000000000003004c7a010000000000000000000000000000000000000003005a7a010000000000000000000000000000000000000003005a7a01000000000000000000000000000000000000000300627a01000000000000000000000000000000000000000300627a010000000000000000000000000000000000000003006a7a010000000000000000000000000000000000000003006a7a010000000000000000000000000000000000000003007a7a010000000000000000000000000000000000000003007a7a010000000000000000000000000000000000000003008a7a010000000000000000000000000000000000000003008c7a01000000000000000000000000000000000000000300907a01000000000000000000000000000000000000000300987a010000000000000000000000000000000000000003009a7a010000000000000000000000000000000000000003009a7a01000000000000000000000000000000000000000300a07a01000000000000000000000000000000000000000300a07a01000000000000000000000000000000000000000300a07a01000000000000000000000000000000000000000300a07a01000000000000000000000000000000000000000300a07a01000000000000000000000000000000000000000300a07a01000000000000000000000000000000000000000300a27a01000000000000000000000000000000000000000300ac7a01000000000000000000000000000000000000000300bc7a01000000000000000000000000000000000000000300c07a01000000000000000000000000000000000000000300ce7a01000000000000000000000000000000000000000300d07a01000000000000000000000000000000000000000300e27a01000000000000000000000000000000000000000300e67a01000000000000000000000000000000000000000300e87a01000000000000000000000000000000000000000300f27a01000000000000000000000000000000000000000300f67a01000000000000000000000000000000000000000300f67a0100000000000000000000000000f62100000000040038bc0100000000000000000000000000002200000000040040bc01000000000000000000000000000a22000002000300f67a01000000000078030000000000000000000000000300f67a01000000000000000000000000000000000000000300f67a01000000000000000000000000000000000000000300f67a01000000000000000000000000000000000000000300f87a01000000000000000000000000000000000000000300f87a01000000000000000000000000000000000000000300f87a010000000000000000000000000000000000000003000a7b010000000000000000000000000000000000000003000e7b010000000000000000000000000000000000000003000e7b01000000000000000000000000000000000000000300107b01000000000000000000000000000000000000000300107b01000000000000000000000000000000000000000300187b01000000000000000000000000000000000000000300187b010000000000000000000000000000000000000003001c7b01000000000000000000000000000000000000000300207b01000000000000000000000000000000000000000300247b01000000000000000000000000000000000000000300247b01000000000000000000000000000000000000000300287b01000000000000000000000000000000000000000300287b010000000000000000000000000000000000000003003a7b010000000000000000000000000000000000000003003a7b010000000000000000000000000000000000000003003e7b010000000000000000000000000000000000000003003e7b01000000000000000000000000000000000000000300407b01000000000000000000000000000000000000000300447b01000000000000000000000000000000000000000300447b01000000000000000000000000000000000000000300487b01000000000000000000000000000000000000000300487b010000000000000000000000000000000000000003004a7b010000000000000000000000000000000000000003004a7b010000000000000000000000000000000000000003004c7b010000000000000000000000000000000000000003004c7b01000000000000000000000000000000000000000300507b01000000000000000000000000000000000000000300507b01000000000000000000000000000000000000000300587b010000000000000000000000000000000000000003005c7b01000000000000000000000000000000000000000300607b01000000000000000000000000000000000000000300607b01000000000000000000000000000000000000000300647b01000000000000000000000000000000000000000300647b01000000000000000000000000000000000000000300687b01000000000000000000000000000000000000000300687b010000000000000000000000000000000000000003006c7b01000000000000000000000000000000000000000300707b01000000000000000000000000000000000000000300707b01000000000000000000000000000000000000000300727b01000000000000000000000000000000000000000300767b010000000000000000000000000000000000000003007a7b010000000000000000000000000000000000000003007a7b010000000000000000000000000000000000000003007e7b01000000000000000000000000000000000000000300827b01000000000000000000000000000000000000000300867b01000000000000000000000000000000000000000300867b01000000000000000000000000000000000000000300887b010000000000000000000000000000000000000003008c7b01000000000000000000000000000000000000000300907b01000000000000000000000000000000000000000300907b01000000000000000000000000000000000000000300927b01000000000000000000000000000000000000000300927b01000000000000000000000000000000000000000300967b01000000000000000000000000000000000000000300967b01000000000000000000000000000000000000000300b47b01000000000000000000000000000000000000000300b47b01000000000000000000000000000000000000000300b87b01000000000000000000000000000000000000000300b87b01000000000000000000000000000000000000000300bc7b01000000000000000000000000000000000000000300c07b01000000000000000000000000000000000000000300c87b01000000000000000000000000000000000000000300cc7b01000000000000000000000000000000000000000300d07b01000000000000000000000000000000000000000300d47b01000000000000000000000000000000000000000300d87b01000000000000000000000000000000000000000300dc7b01000000000000000000000000000000000000000300dc7b01000000000000000000000000000000000000000300e07b01000000000000000000000000000000000000000300e07b01000000000000000000000000000000000000000300e47b01000000000000000000000000000000000000000300e47b01000000000000000000000000000000000000000300e87b01000000000000000000000000000000000000000300ec7b01000000000000000000000000000000000000000300ec7b01000000000000000000000000000000000000000300f27b01000000000000000000000000000000000000000300f67b01000000000000000000000000000000000000000300f87b01000000000000000000000000000000000000000300f87b01000000000000000000000000000000000000000300fe7b01000000000000000000000000000000000000000300fe7b01000000000000000000000000000000000000000300027c01000000000000000000000000000000000000000300027c01000000000000000000000000000000000000000300047c01000000000000000000000000000000000000000300087c01000000000000000000000000000000000000000300087c010000000000000000000000000000000000000003000c7c010000000000000000000000000000000000000003000c7c01000000000000000000000000000000000000000300147c01000000000000000000000000000000000000000300147c01000000000000000000000000000000000000000300187c01000000000000000000000000000000000000000300187c010000000000000000000000000000000000000003001a7c010000000000000000000000000000000000000003001a7c010000000000000000000000000000000000000003001e7c010000000000000000000000000000000000000003001e7c01000000000000000000000000000000000000000300227c01000000000000000000000000000000000000000300227c01000000000000000000000000000000000000000300247c01000000000000000000000000000000000000000300247c01000000000000000000000000000000000000000300267c01000000000000000000000000000000000000000300267c010000000000000000000000000000000000000003002a7c010000000000000000000000000000000000000003002e7c01000000000000000000000000000000000000000300367c01000000000000000000000000000000000000000300367c010000000000000000000000000000000000000003003a7c010000000000000000000000000000000000000003003c7c010000000000000000000000000000000000000003003c7c01000000000000000000000000000000000000000300407c01000000000000000000000000000000000000000300407c01000000000000000000000000000000000000000300447c01000000000000000000000000000000000000000300487c01000000000000000000000000000000000000000300487c010000000000000000000000000000000000000003004a7c010000000000000000000000000000000000000003004a7c01000000000000000000000000000000000000000300527c01000000000000000000000000000000000000000300527c01000000000000000000000000000000000000000300547c01000000000000000000000000000000000000000300547c01000000000000000000000000000000000000000300567c01000000000000000000000000000000000000000300567c010000000000000000000000000000000000000003005a7c010000000000000000000000000000000000000003005a7c01000000000000000000000000000000000000000300607c01000000000000000000000000000000000000000300607c01000000000000000000000000000000000000000300687c01000000000000000000000000000000000000000300687c010000000000000000000000000000000000000003006e7c010000000000000000000000000000000000000003006e7c01000000000000000000000000000000000000000300727c01000000000000000000000000000000000000000300727c01000000000000000000000000000000000000000300747c01000000000000000000000000000000000000000300787c01000000000000000000000000000000000000000300787c010000000000000000000000000000000000000003007a7c010000000000000000000000000000000000000003007a7c01000000000000000000000000000000000000000300827c01000000000000000000000000000000000000000300827c01000000000000000000000000000000000000000300847c01000000000000000000000000000000000000000300847c01000000000000000000000000000000000000000300867c01000000000000000000000000000000000000000300867c01000000000000000000000000000000000000000300887c01000000000000000000000000000000000000000300887c010000000000000000000000000000000000000003008a7c010000000000000000000000000000000000000003008a7c010000000000000000000000000000000000000003008c7c010000000000000000000000000000000000000003008c7c01000000000000000000000000000000000000000300927c01000000000000000000000000000000000000000300967c01000000000000000000000000000000000000000300967c01000000000000000000000000000000000000000300987c01000000000000000000000000000000000000000300987c01000000000000000000000000000000000000000300a07c01000000000000000000000000000000000000000300a07c01000000000000000000000000000000000000000300a27c01000000000000000000000000000000000000000300a27c01000000000000000000000000000000000000000300a47c01000000000000000000000000000000000000000300a47c01000000000000000000000000000000000000000300a67c01000000000000000000000000000000000000000300a67c01000000000000000000000000003922000000000300aa7c01000000000000000000000000004722000000000300b27c01000000000000000000000000000000000000000300c87c01000000000000000000000000000000000000000300ce7c01000000000000000000000000000000000000000300dc7c01000000000000000000000000000000000000000300dc7c01000000000000000000000000000000000000000300e07c01000000000000000000000000000000000000000300e27c01000000000000000000000000000000000000000300e67c01000000000000000000000000000000000000000300e87c01000000000000000000000000000000000000000300e87c01000000000000000000000000000000000000000300ec7c01000000000000000000000000000000000000000300ec7c01000000000000000000000000000000000000000300ee7c01000000000000000000000000000000000000000300ee7c01000000000000000000000000000000000000000300f07c01000000000000000000000000000000000000000300f27c01000000000000000000000000000000000000000300f27c01000000000000000000000000000000000000000300f47c01000000000000000000000000000000000000000300fe7c01000000000000000000000000000000000000000300027d01000000000000000000000000000000000000000300067d01000000000000000000000000000000000000000300067d010000000000000000000000000000000000000003000a7d010000000000000000000000000000000000000003000a7d01000000000000000000000000000000000000000300107d01000000000000000000000000000000000000000300107d01000000000000000000000000000000000000000300127d01000000000000000000000000000000000000000300127d01000000000000000000000000000000000000000300167d01000000000000000000000000000000000000000300187d010000000000000000000000000000000000000003001a7d010000000000000000000000000000000000000003001a7d010000000000000000000000000000000000000003001e7d01000000000000000000000000000000000000000300207d01000000000000000000000000000000000000000300227d01000000000000000000000000000000000000000300227d01000000000000000000000000000000000000000300247d01000000000000000000000000000000000000000300247d01000000000000000000000000000000000000000300287d01000000000000000000000000000000000000000300287d010000000000000000000000000000000000000003002a7d010000000000000000000000000000000000000003002a7d010000000000000000000000000000000000000003002e7d01000000000000000000000000000000000000000300307d01000000000000000000000000000000000000000300307d01000000000000000000000000000000000000000300327d01000000000000000000000000000000000000000300327d01000000000000000000000000000000000000000300347d01000000000000000000000000000000000000000300387d010000000000000000000000000000000000000003003c7d010000000000000000000000000000000000000003003e7d01000000000000000000000000000000000000000300407d01000000000000000000000000000000000000000300427d01000000000000000000000000000000000000000300427d01000000000000000000000000000000000000000300447d01000000000000000000000000000000000000000300447d01000000000000000000000000000000000000000300467d01000000000000000000000000000000000000000300467d010000000000000000000000000000000000000003004a7d010000000000000000000000000000000000000003004a7d010000000000000000000000000000000000000003004e7d01000000000000000000000000000000000000000300507d01000000000000000000000000000000000000000300527d01000000000000000000000000000000000000000300567d01000000000000000000000000000000000000000300567d010000000000000000000000000000000000000003005a7d010000000000000000000000000000000000000003005a7d010000000000000000000000000000000000000003005c7d010000000000000000000000000000000000000003005c7d01000000000000000000000000000000000000000300627d01000000000000000000000000000000000000000300627d01000000000000000000000000000000000000000300667d010000000000000000000000000000000000000003006a7d010000000000000000000000000000000000000003006e7d01000000000000000000000000000000000000000300747d010000000000000000000000000000000000000003007a7d010000000000000000000000000000000000000003007a7d010000000000000000000000000000000000000003007c7d010000000000000000000000000000000000000003007c7d010000000000000000000000000000000000000003007e7d010000000000000000000000000000000000000003007e7d01000000000000000000000000000000000000000300827d01000000000000000000000000000000000000000300847d01000000000000000000000000000000000000000300867d010000000000000000000000000000000000000003008a7d010000000000000000000000000000000000000003008a7d010000000000000000000000000000000000000003008c7d010000000000000000000000000000000000000003008c7d010000000000000000000000000000000000000003008e7d010000000000000000000000000000000000000003008e7d01000000000000000000000000000000000000000300927d01000000000000000000000000000000000000000300927d01000000000000000000000000000000000000000300947d01000000000000000000000000000000000000000300947d01000000000000000000000000000000000000000300987d010000000000000000000000000000000000000003009a7d010000000000000000000000000000000000000003009e7d01000000000000000000000000000000000000000300a07d01000000000000000000000000000000000000000300a07d01000000000000000000000000000000000000000300a47d01000000000000000000000000000000000000000300a47d01000000000000000000000000000000000000000300a67d01000000000000000000000000000000000000000300a67d01000000000000000000000000000000000000000300a87d01000000000000000000000000000000000000000300a87d01000000000000000000000000000000000000000300ac7d01000000000000000000000000000000000000000300ac7d01000000000000000000000000000000000000000300b27d01000000000000000000000000000000000000000300b27d01000000000000000000000000000000000000000300b67d01000000000000000000000000000000000000000300b67d01000000000000000000000000000000000000000300bc7d01000000000000000000000000000000000000000300bc7d01000000000000000000000000000000000000000300e27d01000000000000000000000000000000000000000300e27d01000000000000000000000000000000000000000300e67d01000000000000000000000000000000000000000300ea7d01000000000000000000000000000000000000000300ec7d01000000000000000000000000000000000000000300f27d01000000000000000000000000000000000000000300007e01000000000000000000000000000000000000000300047e01000000000000000000000000000000000000000300047e01000000000000000000000000000000000000000300067e01000000000000000000000000000000000000000300067e01000000000000000000000000000000000000000300087e01000000000000000000000000000000000000000300087e01000000000000000000000000000000000000000300147e01000000000000000000000000000000000000000300147e010000000000000000000000000000000000000003001e7e01000000000000000000000000000000000000000300227e01000000000000000000000000000000000000000300307e01000000000000000000000000000000000000000300307e01000000000000000000000000000000000000000300387e01000000000000000000000000000000000000000300387e010000000000000000000000000000000000000003003c7e010000000000000000000000000000000000000003003c7e01000000000000000000000000000000000000000300407e01000000000000000000000000000000000000000300407e01000000000000000000000000000000000000000300507e01000000000000000000000000000000000000000300527e01000000000000000000000000000000000000000300527e01000000000000000000000000000000000000000300567e01000000000000000000000000000000000000000300567e010000000000000000000000000000000000000003006a7e010000000000000000000000000000000000000003006e7e010000000000000000000000000000000000000003006e7e010000000000000000000000000000000000000003006e7e010000000000000000000000000000000000000003006e7e010000000000000000000000000000000000000003006e7e01000000000000000000000000000000000000000300707e01000000000000000000000000000000000000000300707e01000000000000000000000000000000000000000300727e010000000000000000000000000000000000000003007c7e010000000000000000000000000000000000000003007c7e010000000000000000000000000055220000020003007c7e0100000000007e0100000000000000000000000003007c7e010000000000000000000000000000000000000003007c7e010000000000000000000000000000000000000003007c7e010000000000000000000000000000000000000003007e7e010000000000000000000000000000000000000003008e7e01000000000000000000000000000000000000000300947e01000000000000000000000000000000000000000300947e010000000000000000000000000000000000000003009c7e010000000000000000000000000000000000000003009c7e01000000000000000000000000000000000000000300a07e01000000000000000000000000000000000000000300a07e01000000000000000000000000000000000000000300a87e01000000000000000000000000000000000000000300a87e01000000000000000000000000000000000000000300aa7e01000000000000000000000000000000000000000300ae7e01000000000000000000000000000000000000000300ae7e01000000000000000000000000000000000000000300b27e01000000000000000000000000000000000000000300b67e01000000000000000000000000007c22000000000300d07e01000000000000000000000000000000000000000300d87e01000000000000000000000000000000000000000300d87e01000000000000000000000000000000000000000300da7e01000000000000000000000000000000000000000300dc7e01000000000000000000000000000000000000000300e07e01000000000000000000000000000000000000000300e47e01000000000000000000000000000000000000000300ea7e01000000000000000000000000000000000000000300ea7e01000000000000000000000000000000000000000300ec7e01000000000000000000000000000000000000000300ee7e01000000000000000000000000000000000000000300f27e01000000000000000000000000000000000000000300f67e01000000000000000000000000000000000000000300f87e01000000000000000000000000000000000000000300f87e01000000000000000000000000000000000000000300fc7e01000000000000000000000000000000000000000300fc7e01000000000000000000000000000000000000000300fe7e01000000000000000000000000000000000000000300047f01000000000000000000000000000000000000000300047f010000000000000000000000000000000000000003000a7f010000000000000000000000000000000000000003000a7f01000000000000000000000000000000000000000300147f01000000000000000000000000000000000000000300187f010000000000000000000000000000000000000003001a7f010000000000000000000000000000000000000003001c7f010000000000000000000000000000000000000003001c7f010000000000000000000000000000000000000003001e7f01000000000000000000000000000000000000000300227f010000000000000000000000000000000000000003002a7f010000000000000000000000000000000000000003002a7f01000000000000000000000000000000000000000300307f01000000000000000000000000000000000000000300307f010000000000000000000000000000000000000003003a7f010000000000000000000000000000000000000003003e7f01000000000000000000000000000000000000000300407f01000000000000000000000000000000000000000300427f01000000000000000000000000000000000000000300427f01000000000000000000000000000000000000000300447f01000000000000000000000000000000000000000300487f010000000000000000000000000000000000000003004a7f010000000000000000000000000000000000000003004a7f010000000000000000000000000000000000000003004e7f010000000000000000000000000000000000000003004e7f01000000000000000000000000000000000000000300507f01000000000000000000000000000000000000000300527f01000000000000000000000000000000000000000300567f01000000000000000000000000000000000000000300567f01000000000000000000000000000000000000000300587f01000000000000000000000000000000000000000300587f01000000000000000000000000000000000000000300687f01000000000000000000000000000000000000000300687f010000000000000000000000000000000000000003006c7f010000000000000000000000000000000000000003006c7f01000000000000000000000000000000000000000300707f01000000000000000000000000000000000000000300787f010000000000000000000000000000000000000003008a7f010000000000000000000000000000000000000003008a7f010000000000000000000000000000000000000003008c7f010000000000000000000000000000000000000003008e7f01000000000000000000000000000000000000000300927f01000000000000000000000000000000000000000300967f010000000000000000000000000000000000000003009c7f010000000000000000000000000000000000000003009c7f010000000000000000000000000000000000000003009e7f01000000000000000000000000000000000000000300a27f01000000000000000000000000000000000000000300a67f01000000000000000000000000000000000000000300a67f01000000000000000000000000000000000000000300a87f01000000000000000000000000000000000000000300a87f01000000000000000000000000000000000000000300b27f01000000000000000000000000000000000000000300b27f01000000000000000000000000000000000000000300b67f01000000000000000000000000000000000000000300b67f01000000000000000000000000000000000000000300bc7f01000000000000000000000000000000000000000300bc7f01000000000000000000000000000000000000000300be7f01000000000000000000000000000000000000000300c27f01000000000000000000000000000000000000000300c27f01000000000000000000000000000000000000000300c67f01000000000000000000000000000000000000000300c67f01000000000000000000000000000000000000000300ca7f01000000000000000000000000000000000000000300ca7f01000000000000000000000000000000000000000300ce7f01000000000000000000000000000000000000000300ce7f01000000000000000000000000000000000000000300d27f01000000000000000000000000000000000000000300da7f01000000000000000000000000000000000000000300e07f01000000000000000000000000000000000000000300e67f01000000000000000000000000000000000000000300f67f01000000000000000000000000000000000000000300fa7f01000000000000000000000000000000000000000300fa7f01000000000000000000000000008a22000002000300fa7f01000000000012000000000000000000000000000300fa7f01000000000000000000000000000000000000000300fa7f01000000000000000000000000000000000000000300fa7f01000000000000000000000000000000000000000300fa7f0100000000000000000000000000e42200000000030000800100000000000000000000000000f2220000010001003b050100000000000b0000000000000000000000000003000c80010000000000000000000000000000000000000003000c80010000000000000000000000000000000000000003000c8001000000000000000000000000001e230000020003000c80010000000000120000000000000000000000000003000c80010000000000000000000000000000000000000003000c80010000000000000000000000000000000000000003000c80010000000000000000000000000000000000000003000c8001000000000000000000000000007b2300000000030012800100000000000000000000000000892300000100010046050100000000000e0000000000000000000000000003001e80010000000000000000000000000000000000000003001e80010000000000000000000000000000000000000003001e80010000000000000000000000000000000000000003001e80010000000000000000000000000000000000000003001e80010000000000000000000000000000000000000003001e80010000000000000000000000000000000000000003002080010000000000000000000000000000000000000003002080010000000000000000000000000000000000000003002280010000000000000000000000000000000000000003002c80010000000000000000000000000000000000000003002c80010000000000000000000000000000000000000003002c80010000000000000000000000000000000000000003002c80010000000000000000000000000000000000000003002c80010000000000000000000000000000000000000003002e80010000000000000000000000000000000000000003002e80010000000000000000000000000000000000000003002e80010000000000000000000000000000000000000003003080010000000000000000000000000000000000000003003a80010000000000000000000000000000000000000003003a80010000000000000000000000000000000000000003003a80010000000000000000000000000000000000000003003a80010000000000000000000000000000000000000003003a80010000000000000000000000000000000000000003003a80010000000000000000000000000000000000000003003c80010000000000000000000000000000000000000003003c80010000000000000000000000000000000000000003003e800100000000000000000000000000000000000000030048800100000000000000000000000000000000000000030048800100000000000000000000000000b5230000020003004880010000000000700000000000000000000000000003004880010000000000000000000000000000000000000003004880010000000000000000000000000000000000000003004880010000000000000000000000000000000000000003004a80010000000000000000000000000000000000000003004c80010000000000000000000000000000000000000003004e80010000000000000000000000000000000000000003004e80010000000000000000000000000000000000000003005680010000000000000000000000000000000000000003005680010000000000000000000000000000000000000003005e80010000000000000000000000000000000000000003005e80010000000000000000000000000000000000000003006080010000000000000000000000000000000000000003006080010000000000000000000000000000000000000003006480010000000000000000000000000000000000000003006480010000000000000000000000000000000000000003006c80010000000000000000000000000000000000000003006e80010000000000000000000000000000000000000003006e80010000000000000000000000000000000000000003007680010000000000000000000000000000000000000003007680010000000000000000000000000000000000000003007a80010000000000000000000000000000000000000003007a80010000000000000000000000000000000000000003008480010000000000000000000000000000000000000003008480010000000000000000000000000000000000000003008e80010000000000000000000000000015240000000003008e80010000000000000000000000000023240000010001009c05010000000000020000000000000000000000000003008e8001000000000000000000000000000000000000000300a48001000000000000000000000000000000000000000300a48001000000000000000000000000000000000000000300a68001000000000000000000000000000000000000000300aa8001000000000000000000000000000000000000000300aa8001000000000000000000000000000000000000000300b88001000000000000000000000000000000000000000300b88001000000000000000000000000000000000000000300b88001000000000000000000000000004f2400000000040048bc0100000000000000000000000000592400000000040050bc0100000000000000000000000000632400000000040058bc01000000000000000000000000006d24000002000300b880010000000000bc010000000000000000000000000300b88001000000000000000000000000000000000000000300b88001000000000000000000000000000000000000000300b88001000000000000000000000000000000000000000300ba8001000000000000000000000000000000000000000300d4800100000000000000000000000000d524000000000300de800100000000000000000000000000e324000000000300e6800100000000000000000000000000f124000000000300ee8001000000000000000000000000000000000000000300fe8001000000000000000000000000000000000000000300fe800100000000000000000000000000ff240000000003000681010000000000000000000000000000000000000003001681010000000000000000000000000000000000000003001681010000000000000000000000000000000000000003001a81010000000000000000000000000000000000000003001a81010000000000000000000000000000000000000003002481010000000000000000000000000000000000000003002481010000000000000000000000000000000000000003002881010000000000000000000000000000000000000003003681010000000000000000000000000000000000000003003681010000000000000000000000000000000000000003003e81010000000000000000000000000000000000000003003e81010000000000000000000000000000000000000003004881010000000000000000000000000000000000000003004881010000000000000000000000000000000000000003005081010000000000000000000000000000000000000003005081010000000000000000000000000000000000000003005681010000000000000000000000000000000000000003005681010000000000000000000000000000000000000003005a81010000000000000000000000000000000000000003005c81010000000000000000000000000000000000000003006881010000000000000000000000000000000000000003006a81010000000000000000000000000000000000000003007081010000000000000000000000000000000000000003007081010000000000000000000000000000000000000003007881010000000000000000000000000000000000000003007c81010000000000000000000000000000000000000003007c81010000000000000000000000000000000000000003008a81010000000000000000000000000000000000000003009081010000000000000000000000000000000000000003009481010000000000000000000000000000000000000003009481010000000000000000000000000000000000000003009881010000000000000000000000000000000000000003009881010000000000000000000000000000000000000003009e8101000000000000000000000000000000000000000300a08101000000000000000000000000000000000000000300a08101000000000000000000000000000000000000000300a28101000000000000000000000000000000000000000300a28101000000000000000000000000000000000000000300aa8101000000000000000000000000000000000000000300aa8101000000000000000000000000000000000000000300b48101000000000000000000000000000000000000000300b68101000000000000000000000000000000000000000300b68101000000000000000000000000000000000000000300b88101000000000000000000000000000000000000000300b88101000000000000000000000000000000000000000300c08101000000000000000000000000000000000000000300c08101000000000000000000000000000000000000000300c28101000000000000000000000000000000000000000300c88101000000000000000000000000000000000000000300c88101000000000000000000000000000000000000000300d48101000000000000000000000000000000000000000300d68101000000000000000000000000000000000000000300da8101000000000000000000000000000000000000000300da8101000000000000000000000000000000000000000300de8101000000000000000000000000000000000000000300e28101000000000000000000000000000000000000000300e88101000000000000000000000000000000000000000300e88101000000000000000000000000000000000000000300f48101000000000000000000000000000000000000000300fc8101000000000000000000000000000000000000000300fc8101000000000000000000000000000000000000000300fe81010000000000000000000000000000000000000003000082010000000000000000000000000000000000000003000882010000000000000000000000000000000000000003000882010000000000000000000000000000000000000003000a82010000000000000000000000000000000000000003000a82010000000000000000000000000000000000000003000e82010000000000000000000000000000000000000003000e82010000000000000000000000000000000000000003001282010000000000000000000000000000000000000003001282010000000000000000000000000000000000000003002682010000000000000000000000000000000000000003002c82010000000000000000000000000000000000000003003a8201000000000000000000000000000000000000000300428201000000000000000000000000000000000000000300428201000000000000000000000000000000000000000300468201000000000000000000000000000000000000000300468201000000000000000000000000000000000000000300568201000000000000000000000000000000000000000300708201000000000000000000000000000000000000000300748201000000000000000000000000000000000000000300748201000000000000000000000000000d250000020003007482010000000000b40000000000000000000000000003007482010000000000000000000000000000000000000003007482010000000000000000000000000000000000000003007482010000000000000000000000000000000000000003007682010000000000000000000000000000000000000003007882010000000000000000000000000000000000000003008082010000000000000000000000000000000000000003008282010000000000000000000000000000000000000003008282010000000000000000000000000000000000000003008682010000000000000000000000000000000000000003008682010000000000000000000000000000000000000003008e82010000000000000000000000000000000000000003008e8201000000000000000000000000000000000000000300948201000000000000000000000000000000000000000300948201000000000000000000000000000000000000000300988201000000000000000000000000000000000000000300a08201000000000000000000000000000000000000000300a48201000000000000000000000000000000000000000300b08201000000000000000000000000000000000000000300b08201000000000000000000000000000000000000000300b68201000000000000000000000000000000000000000300b68201000000000000000000000000000000000000000300ba8201000000000000000000000000000000000000000300c28201000000000000000000000000000000000000000300c88201000000000000000000000000000000000000000300d08201000000000000000000000000000000000000000300d48201000000000000000000000000000000000000000300e08201000000000000000000000000000000000000000300e68201000000000000000000000000000000000000000300ee8201000000000000000000000000000000000000000300f48201000000000000000000000000000000000000000300fc82010000000000000000000000000000000000000003000283010000000000000000000000000000000000000003000a83010000000000000000000000000000000000000003000e83010000000000000000000000000000000000000003001883010000000000000000000000000000000000000003001883010000000000000000000000000000000000000003002283010000000000000000000000000000000000000003002483010000000000000000000000000000000000000003002883010000000000000000000000000000000000000003002883010000000000000000000000000040250000020003002883010000000000380000000000000000000000000003002883010000000000000000000000000000000000000003002883010000000000000000000000000000000000000003002883010000000000000000000000000000000000000003002a83010000000000000000000000000000000000000003002a83010000000000000000000000000000000000000003002c8301000000000000000000000000007125000000000300468301000000000000000000000000007f250000010001006806010000000000300000000000000000000000000003005a83010000000000000000000000000000000000000003005c830100000000000000000000000000000000000000030060830100000000000000000000000000000000000000030060830100000000000000000000000000ab2500000200030060830100000000000a0000000000000000000000000003006083010000000000000000000000000000000000000003006083010000000000000000000000000000000000000003006083010000000000000000000000000000000000000003006083010000000000000000000000000000000000000003006a83010000000000000000000000000000000000000003006a83010000000000000000000000000001260000020003006a83010000000000b60000000000000000000000000003006a83010000000000000000000000000000000000000003006a83010000000000000000000000000000000000000003006a83010000000000000000000000000000000000000003006c83010000000000000000000000000000000000000003006c83010000000000000000000000000000000000000003006e83010000000000000000000000000000000000000003007883010000000000000000000000000000000000000003007883010000000000000000000000000000000000000003007a83010000000000000000000000000000000000000003007a83010000000000000000000000000000000000000003007e83010000000000000000000000000000000000000003007e83010000000000000000000000000000000000000003008683010000000000000000000000000000000000000003008683010000000000000000000000000000000000000003008c83010000000000000000000000000000000000000003008c83010000000000000000000000000000000000000003009083010000000000000000000000000000000000000003009883010000000000000000000000000000000000000003009c8301000000000000000000000000000000000000000300a88301000000000000000000000000000000000000000300a88301000000000000000000000000000000000000000300ae8301000000000000000000000000000000000000000300ae8301000000000000000000000000000000000000000300b28301000000000000000000000000000000000000000300ba8301000000000000000000000000000000000000000300c08301000000000000000000000000000000000000000300c88301000000000000000000000000000000000000000300cc8301000000000000000000000000000000000000000300d88301000000000000000000000000000000000000000300de8301000000000000000000000000000000000000000300e68301000000000000000000000000000000000000000300ec8301000000000000000000000000000000000000000300f48301000000000000000000000000000000000000000300fa83010000000000000000000000000000000000000003000284010000000000000000000000000000000000000003000684010000000000000000000000000000000000000003001084010000000000000000000000000000000000000003001084010000000000000000000000000000000000000003001a84010000000000000000000000000000000000000003001a84010000000000000000000000000000000000000003001c840100000000000000000000000000000000000000030020840100000000000000000000000000000000000000030020840100000000000000000000000000592600000200030020840100000000003a00000000000000000000000000030020840100000000000000000000000000000000000000030020840100000000000000000000000000000000000000030020840100000000000000000000000000000000000000030022840100000000000000000000000000000000000000030022840100000000000000000000000000000000000000030024840100000000000000000000000000af260000000003004084010000000000000000000000000000000000000003004084010000000000000000000000000000000000000003004084010000000000000000000000000000000000000003005484010000000000000000000000000000000000000003005484010000000000000000000000000000000000000003005684010000000000000000000000000000000000000003005a84010000000000000000000000000000000000000003005a840100000000000000000000000000bd260000020003005a84010000000000200100000000000000000000000003005a84010000000000000000000000000000000000000003005a84010000000000000000000000000000000000000003005a84010000000000000000000000000000000000000003005c84010000000000000000000000000000000000000003006a84010000000000000000000000000000000000000003006c84010000000000000000000000000000000000000003007084010000000000000000000000000000000000000003007084010000000000000000000000000000000000000003007284010000000000000000000000000000000000000003007284010000000000000000000000000000000000000003007a84010000000000000000000000000000000000000003007e84010000000000000000000000000000000000000003007e84010000000000000000000000000000000000000003008284010000000000000000000000000000000000000003008284010000000000000000000000000000000000000003008684010000000000000000000000000000000000000003008684010000000000000000000000000000000000000003008a84010000000000000000000000000000000000000003008a84010000000000000000000000000000000000000003008e84010000000000000000000000000000000000000003008e840100000000000000000000000000000000000000030090840100000000000000000000000000000000000000030094840100000000000000000000000000f926000000000300988401000000000000000000000000000727000001000100960501000000000002000000000000000000000000000300988401000000000000000000000000000000000000000300a28401000000000000000000000000000000000000000300a68401000000000000000000000000000000000000000300a68401000000000000000000000000003327000000000300b08401000000000000000000000000004127000001000100980501000000000002000000000000000000000000000300bc8401000000000000000000000000000000000000000300bc8401000000000000000000000000000000000000000300be8401000000000000000000000000006d27000000000300c48401000000000000000000000000007b270000010001009a0501000000000001000000000000000000000000000300cc8401000000000000000000000000000000000000000300cc8401000000000000000000000000000000000000000300d68401000000000000000000000000000000000000000300d68401000000000000000000000000000000000000000300d88401000000000000000000000000000000000000000300d88401000000000000000000000000000000000000000300dc8401000000000000000000000000000000000000000300dc8401000000000000000000000000000000000000000300de8401000000000000000000000000000000000000000300de8401000000000000000000000000000000000000000300ea8401000000000000000000000000000000000000000300ea8401000000000000000000000000000000000000000300ee8401000000000000000000000000000000000000000300ee8401000000000000000000000000000000000000000300f08401000000000000000000000000000000000000000300f48401000000000000000000000000000000000000000300f48401000000000000000000000000000000000000000300fc8401000000000000000000000000000000000000000300fc84010000000000000000000000000000000000000003000685010000000000000000000000000000000000000003000685010000000000000000000000000000000000000003000a85010000000000000000000000000000000000000003000e85010000000000000000000000000000000000000003001685010000000000000000000000000000000000000003001e850100000000000000000000000000000000000000030032850100000000000000000000000000000000000000030032850100000000000000000000000000000000000000030036850100000000000000000000000000a72700000000030036850100000000000000000000000000b52700000100010058050100000000003000000000000000000000000000030036850100000000000000000000000000000000000000030040850100000000000000000000000000000000000000030040850100000000000000000000000000000000000000030048850100000000000000000000000000000000000000030048850100000000000000000000000000e1270000000003004e850100000000000000000000000000ef270000010001009405010000000000020000000000000000000000000003005a85010000000000000000000000000000000000000003005a85010000000000000000000000000000000000000003005c85010000000000000000000000000000000000000003005c85010000000000000000000000000000000000000003006085010000000000000000000000000000000000000003006685010000000000000000000000000000000000000003007685010000000000000000000000000000000000000003007a85010000000000000000000000000000000000000003007a85010000000000000000000000000000000000000003007a85010000000000000000000000000000000000000003007a85010000000000000000000000000000000000000003007a85010000000000000000000000000000000000000003007c85010000000000000000000000000000000000000003008485010000000000000000000000000000000000000003008685010000000000000000000000000000000000000003008685010000000000000000000000000000000000000003009285010000000000000000000000000000000000000003009285010000000000000000000000000000000000000003009e85010000000000000000000000000000000000000003009e8501000000000000000000000000000000000000000300ac8501000000000000000000000000000000000000000300ac8501000000000000000000000000000000000000000300ae8501000000000000000000000000000000000000000300b28501000000000000000000000000000000000000000300b48501000000000000000000000000000000000000000300b68501000000000000000000000000000000000000000300b68501000000000000000000000000000000000000000300b88501000000000000000000000000000000000000000300b88501000000000000000000000000000000000000000300c28501000000000000000000000000000000000000000300c48501000000000000000000000000000000000000000300cc8501000000000000000000000000000000000000000300cc8501000000000000000000000000000000000000000300d28501000000000000000000000000000000000000000300d28501000000000000000000000000000000000000000300d48501000000000000000000000000000000000000000300d48501000000000000000000000000001b28000000000300da85010000000000000000000000000029280000010001009b0501000000000001000000000000000000000000000300e88501000000000000000000000000000000000000000300e88501000000000000000000000000000000000000000300ea8501000000000000000000000000000000000000000300ea8501000000000000000000000000005528000000000300f085010000000000000000000000000063280000010001003a05010000000000010000000000000000000000000003000086010000000000000000000000000000000000000003000086010000000000000000000000000000000000000003000486010000000000000000000000000000000000000003000486010000000000000000000000000000000000000003000e8601000000000000000000000000000000000000000300128601000000000000000000000000000000000000000300128601000000000000000000000000000000000000000300128601000000000000000000000000000000000000000300128601000000000000000000000000000000000000000300128601000000000000000000000000000000000000000300148601000000000000000000000000000000000000000300148601000000000000000000000000000000000000000300168601000000000000000000000000000000000000000300208601000000000000000000000000000000000000000300208601000000000000000000000000008f2800000200030020860100000000001600000000000000000000000000030020860100000000000000000000000000000000000000030020860100000000000000000000000000d72800000000030020860100000000000000000000000000000000000000030020860100000000000000000000000000e5280000010001009806010000000000020000000000000000000000000003002086010000000000000000000000000000000000000003003686010000000000000000000000000000000000000003003686010000000000000000000000000000000000000003003686010000000000000000000000000011290000020003003686010000000000a20000000000000000000000000003003686010000000000000000000000000000000000000003003686010000000000000000000000000000000000000003003686010000000000000000000000000000000000000003003886010000000000000000000000000000000000000003003e8601000000000000000000000000000000000000000300408601000000000000000000000000000000000000000300408601000000000000000000000000000000000000000300428601000000000000000000000000000000000000000300428601000000000000000000000000000000000000000300448601000000000000000000000000000000000000000300448601000000000000000000000000007229000000000300488601000000000000000000000000008029000001000100c0060100000000001100000000000000000000000000030054860100000000000000000000000000000000000000030054860100000000000000000000000000000000000000030060860100000000000000000000000000ac2900000000030060860100000000000000000000000000ba29000001000100a006010000000000200000000000000000000000000003006086010000000000000000000000000000000000000003007486010000000000000000000000000000000000000003007486010000000000000000000000000000000000000003007686010000000000000000000000000000000000000003007a86010000000000000000000000000000000000000003007c86010000000000000000000000000000000000000003007e86010000000000000000000000000000000000000003007e86010000000000000000000000000000000000000003008086010000000000000000000000000000000000000003008086010000000000000000000000000000000000000003008a86010000000000000000000000000000000000000003008c86010000000000000000000000000000000000000003009486010000000000000000000000000000000000000003009486010000000000000000000000000000000000000003009a86010000000000000000000000000000000000000003009a86010000000000000000000000000000000000000003009c86010000000000000000000000000000000000000003009c860100000000000000000000000000e629000000000300a28601000000000000000000000000000000000000000300b08601000000000000000000000000000000000000000300b08601000000000000000000000000000000000000000300b28601000000000000000000000000000000000000000300b2860100000000000000000000000000f429000000000300b88601000000000000000000000000000000000000000300c88601000000000000000000000000000000000000000300c88601000000000000000000000000000000000000000300cc8601000000000000000000000000000000000000000300cc8601000000000000000000000000000000000000000300d48601000000000000000000000000000000000000000300d88601000000000000000000000000000000000000000300d8860100000000000000000000000000022a000002000300d88601000000000070000000000000000000000000000300d88601000000000000000000000000000000000000000300d88601000000000000000000000000000000000000000300d88601000000000000000000000000000000000000000300da8601000000000000000000000000000000000000000300dc8601000000000000000000000000000000000000000300de8601000000000000000000000000000000000000000300de8601000000000000000000000000000000000000000300e68601000000000000000000000000000000000000000300e68601000000000000000000000000000000000000000300ee8601000000000000000000000000000000000000000300ee8601000000000000000000000000000000000000000300f08601000000000000000000000000000000000000000300f08601000000000000000000000000000000000000000300f48601000000000000000000000000000000000000000300f48601000000000000000000000000000000000000000300fc8601000000000000000000000000000000000000000300fe8601000000000000000000000000000000000000000300fe86010000000000000000000000000000000000000003000687010000000000000000000000000000000000000003000687010000000000000000000000000000000000000003000a87010000000000000000000000000000000000000003000a87010000000000000000000000000000000000000003001487010000000000000000000000000000000000000003001487010000000000000000000000000000000000000003001e870100000000000000000000000000622a0000000003001e87010000000000000000000000000000000000000003001e87010000000000000000000000000000000000000003003487010000000000000000000000000000000000000003003487010000000000000000000000000000000000000003003687010000000000000000000000000000000000000003003a87010000000000000000000000000000000000000003003a870100000000000000000000000000000000000000030048870100000000000000000000000000000000000000030048870100000000000000000000000000000000000000030048870100000000000000000000000000702a0000020003004887010000000000520000000000000000000000000003004887010000000000000000000000000000000000000003004a8701000000000000000000000000000000000000000300548701000000000000000000000000001c2b0000020003009a870100000000007e0000000000000000000000000003009a87010000000000000000000000000000000000000003009a87010000000000000000000000000000000000000003009c8701000000000000000000000000000000000000000300a287010000000000000000000000000000000000000003001888010000000000000000000000000000000000000003001888010000000000000000000000000000000000000003001a880100000000000000000000000000000000000000030022880100000000000000000000000000762b000002000300b691010000000000080000000000000000000000000003007a880100000000000000000000000000852b0000020003007a88010000000000300000000000000000000000000003007a8801000000000000000000000000000000000000000300aa8801000000000000000000000000000000000000000300aa8801000000000000000000000000000000000000000300ac8801000000000000000000000000000000000000000300b0880100000000000000000000000000cd2b000002000300be9101000000000008000000000000000000000000000300f8880100000000000000000000000000e12b000002000300f88801000000000068000000000000000000000000000300f88801000000000000000000000000000000000000000300fa880100000000000000000000000000000000000000030004890100000000000000000000000000222c00000200030060890100000000007e000000000000000000000000000300608901000000000000000000000000000000000000000300608901000000000000000000000000000000000000000300628901000000000000000000000000000000000000000300688901000000000000000000000000007c2c000002000300de8901000000000052000000000000000000000000000300de8901000000000000000000000000000000000000000300de8901000000000000000000000000000000000000000300e08901000000000000000000000000000000000000000300e68901000000000000000000000000000000000000000300308a01000000000000000000000000000000000000000300308a01000000000000000000000000000000000000000300328a01000000000000000000000000000000000000000300368a01000000000000000000000000000000000000000300868a0100000000000000000000000000af2c000002000300868a01000000000082010000000000000000000000000300868a01000000000000000000000000000000000000000300888a01000000000000000000000000000000000000000300968a0100000000000000000000000000e02c000000000300688b0100000000000000000000000000ee2c000001000100a0070100000000001c00000000000000f82c000000000300728b0100000000000000000000000000062d0000000003007c8b0100000000000000000000000000142d000000000300908b0100000000000000000000000000222d000000000300988b0100000000000000000000000000302d000001000100f80601000000000020000000000000005a2d000000000300a68b0100000000000000000000000000682d00000100010006080100000000002f00000000000000932d000000000300b48b0100000000000000000000000000a12d00000100010035080100000000003200000000000000cc2d000000000300ce8b0100000000000000000000000000da2d000000000300d68b0100000000000000000000000000e82d00000100010080070100000000002000000000000000122e000000000300f08b0100000000000000000000000000202e000001000100bc070100000000001c000000000000004b2e000000000300fa8b0100000000000000000000000000592e000001000100d8070100000000002e000000000000000000000000000300088c0100000000000000000000000000842e000002000300088c01000000000028000000000000000000000000000300088c0100000000000000000000000000df2e0000000003000e8c0100000000000000000000000000ed2e000001000100280a0100000000005000000000000000572f000000000300188c0100000000000000000000000000652f000001000100780a01000000000050000000000000000000000000000300308c0100000000000000000000000000d32f000002000300308c01000000000062000000000000000000000000000300308c01000000000000000000000000000000000000000300328c01000000000000000000000000000c30000000000300528c01000000000000000000000000001a300000000003005e8c01000000000000000000000000002830000001000100180701000000000018000000000000005230000000000300668c01000000000000000000000000006030000001000100300701000000000020000000000000008a300000000003007c8c01000000000000000000000000009830000001000100670801000000000026000000000000000000000000000300928c0100000000000000000000000000c330000002000300928c01000000000068000000000000000000000000000300928c01000000000000000000000000000000000000000300948c01000000000000000000000000000000000000000300988c01000000000000000000000000000231000000000300c48c01000000000000000000000000001031000000000300cc8c01000000000000000000000000001e31000000000300e68c01000000000000000000000000002c310000010001008d080100000000000d000000000000000000000000000300fa8c01000000000000000000000000000000000000000300fa8c01000000000000000000000000000000000000000300fc8c01000000000000000000000000000000000000000300008d01000000000000000000000000005731000000000300388d010000000000000000000000000000000000000003004e8d010000000000000000000000000000000000000003004e8d01000000000000000000000000000000000000000300508d01000000000000000000000000000000000000000300628d01000000000000000000000000006531000000000300e88d01000000000000000000000000007331000000000300768e01000000000000000000000000008131000000000300808e01000000000000000000000000008f310000010001009a080100000000000e00000000000000ba310000000003008c8e0100000000000000000000000000c831000000000300968e0100000000000000000000000000d631000000000300a08e0100000000000000000000000000e431000000000300aa8e0100000000000000000000000000f231000000000300b48e01000000000000000000000000000000000000000300ca8e01000000000000000000000000000000000000000300ca8e01000000000000000000000000000000000000000300cc8e01000000000000000000000000000000000000000300d28e010000000000000000000000000000320000000003000c8f01000000000000000000000000000e32000000000300148f01000000000000000000000000001c320000000003002e8f01000000000000000000000000002a32000001000100a8080100000000000e000000000000000000000000000300428f01000000000000000000000000000000000000000300428f01000000000000000000000000000000000000000300448f010000000000000000000000000000000000000003004a8f010000000000000000000000000055320000000003008a8f01000000000000000000000000006332000000000300928f01000000000000000000000000007132000000000300ac8f01000000000000000000000000007f32000001000100b6080100000000000d000000000000000000000000000300c08f01000000000000000000000000000000000000000300c08f01000000000000000000000000000000000000000300c28f01000000000000000000000000000000000000000300ca8f0100000000000000000000000000aa320000000003002c900100000000000000000000000000b83200000000030034900100000000000000000000000000c6320000000003004e900100000000000000000000000000d432000001000100c3080100000000001200000000000000000000000000030062900100000000000000000000000000ff3200000200030062900100000000007a0000000000000000000000000003006290010000000000000000000000000000000000000003006490010000000000000000000000000000000000000003006a9001000000000000000000000000006333000000000300ba9001000000000000000000000000000000000000000300dc9001000000000000000000000000000000000000000300dc9001000000000000000000000000000000000000000300de9001000000000000000000000000000000000000000300ea9001000000000000000000000000007133000000000300449101000000000000000000000000007f33000001000100d8080100000000002000000000000000000000000000030096910100000000000000000000000000aa33000002000300969101000000000010000000000000000000000000000300969101000000000000000000000000000000000000000300a69101000000000000000000000000000000000000000300a69101000000000000000000000000000000000000000300ae9101000000000000000000000000000000000000000300ae9101000000000000000000000000000000000000000300b69101000000000000000000000000000000000000000300b69101000000000000000000000000000000000000000300be9101000000000000000000000000000000000000000300be9101000000000000000000000000000000000000000300c69101000000000000000000000000000000000000000300c69101000000000000000000000000000000000000000300d09101000000000000000000000000000000000000000300d09101000000000000000000000000000000000000000300d29101000000000000000000000000000000000000000300da910100000000000000000000000000fb330000000003002492010000000000000000000000000000000000000003004292010000000000000000000000000009340000020003004292010000000000ca020000000000000000000000000300429201000000000000000000000000000000000000000300449201000000000000000000000000000000000000000300549201000000000000000000000000009334000000000300ce940100000000000000000000000000a134000000000300e2940100000000000000000000000000af34000000000300ec940100000000000000000000000000bd34000000000300f494010000000000000000000000000000000000000003000c95010000000000000000000000000000000000000003000c950100000000000000000000000000cb340000000003000e950100000000000000000000000000d93400000000010088010100000000000000000000000000e4340000000003001e950100000000000000000000000000ee3400000000030020950100000000000000000000000000f834000000000300229501000000000000000000000000000235000000000300269501000000000000000000000000000c350000000003002a95010000000000000000000000000000000000000003003495010000000000000000000000000000000000000003003495010000000000000000000000000000000000000003003695010000000000000000000000000000000000000003004695010000000000000000000000000000000000000003009896010000000000000000000000000000000000000003009896010000000000000000000000000000000000000003009c9601000000000000000000000000000000000000000300c09601000000000000000000000000001635000000000300209a01000000000000000000000000002435000000000300a29b0100000000000000000000000000323500000100010030040100000000001c000000000000003b35000000000300ac9b01000000000000000000000000004935000000000300b69b01000000000000000000000000005735000000000300c09b01000000000000000000000000006535000000000300ca9b01000000000000000000000000007335000000000300de9b01000000000000000000000000008135000000000300e69b01000000000000000000000000008f350000010001009009010000000000200000000000000000000000000003001e9c010000000000000000000000000000000000000003001e9c01000000000000000000000000000000000000000300209c01000000000000000000000000000000000000000300369c0100000000000000000000000000ba35000000000300f49e0100000000000000000000000000c835000000000300089f0100000000000000000000000000d635000001000100d0090100000000002b000000000000000236000000000300169f010000000000000000000000000010360000000003001e9f01000000000000000000000000000000000000000300369f01000000000000000000000000000000000000000300369f01000000000000000000000000000000000000000300389f010000000000000000000000000000000000000003003e9f01000000000000000000000000000000000000000300c89f01000000000000000000000000000000000000000300c89f01000000000000000000000000000000000000000300ca9f01000000000000000000000000000000000000000300e49f01000000000000000000000000001e360000000003001ca301000000000000000000000000002c3600000000030030a301000000000000000000000000003a3600000000030038a30100000000000000000000000000483600000000030050a301000000000000000000000000005636000001000100fb090100000000002900000000000000000000000000030068a30100000000000000000000000000000000000000030068a3010000000000000000000000000000000000000003006aa30100000000000000000000000000000000000000030076a301000000000000000000000000008236000000000300c8a401000000000000000000000000000000000000000300eea40100000000000000000000000000903600000100060018bd0100000000000010080000000000bb3600000100060018cd0900000000000010000000000000ec360000010001007c0301000000000023000000000000001737000001000100b00301000000000033000000000000004237000001000100f8080100000000000a000000000000006d3700000100010002090100000000000a0000000000000098370000010001000c090100000000000b00000000000000c33700000100010017090100000000000600000000000000ee370000010001001d09010000000000060000000000000019380000010001002309010000000000090000000000000044380000010001002c0901000000000006000000000000000000000000000800000000000000000000000000000000000000000000000b006f2900000000000000000000000000000000000000000b00114300000000000000000000000000006f38000000000f00000000000000000000000000000000000000000000000b00051200000000000000000000000000000000000000000a00700e00000000000000000000000000000000000000000b001e2d00000000000000000000000000000000000000000b00000000000000000000000000000000000000000000000b00c44b00000000000000000000000000000000000000000b00783500000000000000000000000000000000000000000b00463c00000000000000000000000000000000000000000b001d0e00000000000000000000000000000000000000000800740000000000000000000000000000000000000000000b00f91500000000000000000000000000008338000000000f00880000000000000000000000000000000000000000000a00a00e00000000000000000000000000000000000000000b00da1800000000000000000000000000000000000000000b001f0500000000000000000000000000000000000000000b007d0c00000000000000000000000000000000000000000b002f1600000000000000000000000000000000000000000b00f03200000000000000000000000000000000000000000b002b0c00000000000000000000000000000000000000000b005c3c00000000000000000000000000000000000000000b00ab3000000000000000000000000000000000000000000b00fa3500000000000000000000000000000000000000000b00712300000000000000000000000000000000000000000b00942800000000000000000000000000000000000000000b00c52100000000000000000000000000000000000000000b00e52a00000000000000000000000000000000000000000b00194600000000000000000000000000000000000000000b006b3800000000000000000000000000000000000000000b00833700000000000000000000000000000000000000000b00c50b00000000000000000000000000000000000000000b00f90300000000000000000000000000000000000000000b00ad0c00000000000000000000000000000000000000000b005f3f00000000000000000000000000000000000000000b00c43000000000000000000000000000000000000000000b002c1700000000000000000000000000000000000000000b004d0b00000000000000000000000000000000000000000b00e93400000000000000000000000000000000000000000b00a60000000000000000000000000000000000000000000b00c14600000000000000000000000000000000000000000b00d71200000000000000000000000000000000000000000b00084100000000000000000000000000000000000000000b006c4500000000000000000000000000000000000000000b002b0500000000000000000000000000000000000000000b00060800000000000000000000000000000000000000000b00cc0000000000000000000000000000000000000000000b00052800000000000000000000000000000000000000000b00a73000000000000000000000000000000000000000000b00351200000000000000000000000000000000000000000b00a43100000000000000000000000000000000000000000b00454800000000000000000000000000000000000000000b004e2700000000000000000000000000000000000000000b002c3e00000000000000000000000000000000000000000b00101300000000000000000000000000000000000000000b00104600000000000000000000000000000000000000000b00403b00000000000000000000000000000000000000000b009c4800000000000000000000000000000000000000000b00632e00000000000000000000000000000000000000000b009b1500000000000000000000000000000000000000000b008a3500000000000000000000000000000000000000000a00000000000000000000000000000000000000000000000a00400000000000000000000000000000000000000000000a00700000000000000000000000000000000000000000000a00a00000000000000000000000000000000000000000000b00a30b00000000000000000000000000000000000000000b00412b00000000000000000000000000000000000000000b00713b00000000000000000000000000000000000000000b00be2d00000000000000000000000000000000000000000b00482900000000000000000000000000000000000000000b00242900000000000000000000000000000000000000000b00db1300000000000000000000000000000000000000000b00b11b00000000000000000000000000000000000000000b003c4400000000000000000000000000000000000000000b000d4700000000000000000000000000000000000000000b00ce3800000000000000000000000000000000000000000b00501400000000000000000000000000000000000000000b00032e00000000000000000000000000000000000000000a00200900000000000000000000000000000000000000000a00500900000000000000000000000000000000000000000a00800900000000000000000000000000000000000000000a00b00900000000000000000000000000000000000000000a00e00900000000000000000000000000000000000000000b00650700000000000000000000000000000000000000000b00873200000000000000000000000000000000000000000b006f0700000000000000000000000000000000000000000b001f0300000000000000000000000000000000000000000a00800d00000000000000000000000000000000000000000a00b00d00000000000000000000000000000000000000000a00e00d00000000000000000000000000000000000000000a00100e00000000000000000000000000000000000000000a00400e00000000000000000000000000000000000000000b001f4a00000000000000000000000000000000000000000b00370a00000000000000000000000000000000000000000b006c0a00000000000000000000000000000000000000000b007f0300000000000000000000000000000000000000000b00672e00000000000000000000000000000000000000000b00114900000000000000000000000000000000000000000b00f44000000000000000000000000000000000000000000b00b90c00000000000000000000000000000000000000000b00230500000000000000000000000000000000000000000b00890200000000000000000000000000000000000000000b00e03100000000000000000000000000000000000000000a00d00000000000000000000000000000000000000000000a00100100000000000000000000000000000000000000000a00400100000000000000000000000000000000000000000a00700100000000000000000000000000000000000000000a00a00100000000000000000000000000000000000000000a00d00100000000000000000000000000000000000000000a00000200000000000000000000000000000000000000000a00300200000000000000000000000000000000000000000a00800200000000000000000000000000000000000000000b00c04700000000000000000000000000000000000000000b00f92d00000000000000000000000000000000000000000a00b00200000000000000000000000000000000000000000a00e00200000000000000000000000000000000000000000a00100300000000000000000000000000000000000000000a00400300000000000000000000000000000000000000000a00700300000000000000000000000000000000000000000a00a00300000000000000000000000000000000000000000a00d00300000000000000000000000000000000000000000a00000400000000000000000000000000000000000000000a00300400000000000000000000000000000000000000000a00800400000000000000000000000000000000000000000a00b00400000000000000000000000000000000000000000a00000500000000000000000000000000000000000000000a00300500000000000000000000000000000000000000000a00800500000000000000000000000000000000000000000a00b00500000000000000000000000000000000000000000a00f00500000000000000000000000000000000000000000a00600600000000000000000000000000000000000000000a00b00600000000000000000000000000000000000000000a00f00600000000000000000000000000000000000000000a00200700000000000000000000000000000000000000000a00500700000000000000000000000000000000000000000b003c3800000000000000000000000000000000000000000b00ae2d00000000000000000000000000000000000000000b00371700000000000000000000000000000000000000000b00372b00000000000000000000000000000000000000000b00263100000000000000000000000000000000000000000b00172900000000000000000000000000000000000000000b001a2700000000000000000000000000000000000000000b00431c00000000000000000000000000000000000000000b001f0700000000000000000000000000000000000000000b00572300000000000000000000000000000000000000000b001e1a00000000000000000000000000000000000000000b00f81600000000000000000000000000000000000000000b00fb2e00000000000000000000000000000000000000000b00012f00000000000000000000000000000000000000000b00cf4900000000000000000000000000000000000000000b00d81900000000000000000000000000000000000000000b00fa0800000000000000000000000000000000000000000b008b4900000000000000000000000000000000000000000b001b0f00000000000000000000000000000000000000000b001f0900000000000000000000000000000000000000000b00453900000000000000000000000000000000000000000a00800700000000000000000000000000000000000000000a00b00700000000000000000000000000000000000000000a00e00700000000000000000000000000000000000000000a00100800000000000000000000000000000000000000000a00400800000000000000000000000000000000000000000a00700800000000000000000000000000000000000000000a00a00800000000000000000000000000000000000000000a00e00800000000000000000000000000000000000000000b00f10100000000000000000000000000000000000000000b00d53c00000000000000000000000000000000000000000b00bd3800000000000000000000000000000000000000000b00ec3700000000000000000000000000000000000000000b00923500000000000000000000000000000000000000000a00100a00000000000000000000000000000000000000000a00400a00000000000000000000000000000000000000000a00700a00000000000000000000000000000000000000000a00a00a00000000000000000000000000000000000000000a00d00a00000000000000000000000000000000000000000a00000b00000000000000000000000000000000000000000b00623d00000000000000000000000000000000000000000b00f64400000000000000000000000000000000000000000b00920400000000000000000000000000000000000000000b00d11900000000000000000000000000000000000000000b00fc2200000000000000000000000000000000000000000b003d2900000000000000000000000000000000000000000b008f4900000000000000000000000000000000000000000b00ae4600000000000000000000000000000000000000000b00bd0900000000000000000000000000000000000000000a00b00b00000000000000000000000000000000000000000a00e00b00000000000000000000000000000000000000000a00100c00000000000000000000000000000000000000000a00400c00000000000000000000000000000000000000000a00700c00000000000000000000000000000000000000000a00b00c00000000000000000000000000000000000000000b00bd1c00000000000000000000000000000000000000000b00b54700000000000000000000000000000000000000000b00821c00000000000000000000000000000000000000000b00b92d00000000000000000000000000000000000000000b00f10800000000000000000000000000000000000000000b001f3500000000000000000000000000000000000000000b00693100000000000000000000000000000000000000000b00ec2200000000000000000000000000000000000000000b00e82f00000000000000000000000000000000000000000a00300b00000000000000000000000000000000000000000b004d1800000000000000000000000000000000000000000b00ee2f00000000000000000000000000000000000000000b00c54400000000000000000000000000000000000000000b00994b00000000000000000000000000000000000000000b00ef4700000000000000000000000000000000000000000b00284200000000000000000000000000000000000000000b00534200000000000000000000000000000000000000000a00700b00000000000000000000000000000000000000000b00963700000000000000000000000000000000000000000b00780900000000000000000000000000000000000000000b00b40f00000000000000000000000000000000000000000b00210c00000000000000000000000000000000000000000b005f3000000000000000000000000000000000000000000b00ff0f00000000000000000000000000000000000000000b008c3900000000000000000000000000000000000000000b00164a00000000000000000000000000000000000000000b00954800000000000000000000000000000000000000000b00820900000000000000000000000000000000000000000b00fd4b00000000000000000000000000000000000000000b00903900000000000000000000000000000000000000000b00f90900000000000000000000000000000000000000000b00681000000000000000000000000000000000000000000b00b13100000000000000000000000000000000000000000b00fa1c00000000000000000000000000000000000000000b00792300000000000000000000000000000000000000000b007a3300000000000000000000000000000000000000000b00564500000000000000000000000000000000000000000b00c63a00000000000000000000000000000000000000000b00c10100000000000000000000000000000000000000000b006b2a00000000000000000000000000000000000000000b00274100000000000000000000000000000000000000000b00b34a00000000000000000000000000000000000000000b000b3e00000000000000000000000000000000000000000b00f91a00000000000000000000000000000000000000000b00b73c00000000000000000000000000000000000000000b004c3600000000000000000000000000000000000000000b00120000000000000000000000000000000000000000000b00fd1900000000000000000000000000000000000000000b002b2d00000000000000000000000000000000000000000b00514900000000000000000000000000000000000000000b00f53100000000000000000000000000000000000000000b00d52100000000000000000000000000000000000000000b00e52100000000000000000000000000000000000000000b005f3400000000000000000000000000000000000000000b00a94a00000000000000000000000000000000000000000b00033700000000000000000000000000000000000000000b00c20a00000000000000000000000000000000000000000b00b03a00000000000000000000000000000000000000000b009b0b00000000000000000000000000000000000000000b00731b00000000000000000000000000000000000000000b00dd4100000000000000000000000000000000000000000b00641100000000000000000000000000000000000000000b002a1a00000000000000000000000000000000000000000b00a91a00000000000000000000000000000000000000000b00f62700000000000000000000000000000000000000000b00f14300000000000000000000000000000000000000000b00e24600000000000000000000000000000000000000000b00852500000000000000000000000000000000000000000b00ac3d00000000000000000000000000000000000000000b00b30500000000000000000000000000000000000000000b00c33d00000000000000000000000000000000000000000b00434100000000000000000000000000000000000000000b00b00800000000000000000000000000000000000000000b00342800000000000000000000000000000000000000000b00802800000000000000000000000000000000000000000b00f53700000000000000000000000000000000000000000b009f3a00000000000000000000000000000000000000000b00531900000000000000000000000000000000000000000b00ab1100000000000000000000000000000000000000000b00974100000000000000000000000000000000000000000b00432f00000000000000000000000000000000000000000b001f2600000000000000000000000000000000000000000b00280900000000000000000000000000000000000000000b00a90d00000000000000000000000000000000000000000b00ca1700000000000000000000000000000000000000000b004c0400000000000000000000000000000000000000000b00a91900000000000000000000000000000000000000000b000f0700000000000000000000000000000000000000000b00ab4200000000000000000000000000000000000000000b007a3900000000000000000000000000000000000000000b00b40300000000000000000000000000000000000000000b004a0500000000000000000000000000000000000000000b00ed3100000000000000000000000000000000000000000b00753400000000000000000000000000000000000000000b00f02800000000000000000000000000000000000000000b00400d00000000000000000000000000000000000000000b00d91100000000000000000000000000000000000000000b00353e00000000000000000000000000000000000000000b00123100000000000000000000000000000000000000000b008d3700000000000000000000000000000000000000000b00fa0100000000000000000000000000000000000000000b00364600000000000000000000000000000000000000000b00542f00000000000000000000000000000000000000000b006c1700000000000000000000000000000000000000000b00c31400000000000000000000000000000000000000000b00ec0c00000000000000000000000000000000000000000b00594900000000000000000000000000000000000000000b005a1400000000000000000000000000000000000000000b00983b00000000000000000000000000000000000000000b00b71b00000000000000000000000000000000000000000b00573d00000000000000000000000000000000000000000b00b22d00000000000000000000000000000000000000000b00d81700000000000000000000000000000000000000000b00a63b00000000000000000000000000000000000000000b00de3b00000000000000000000000000000000000000000b00744700000000000000000000000000000000000000000b00341c00000000000000000000000000000000000000000b00760f00000000000000000000000000000000000000000b00a93e00000000000000000000000000000000000000000b00242d00000000000000000000000000000000000000000b00b02900000000000000000000000000000000000000000b00494300000000000000000000000000000000000000000b00381200000000000000000000000000000000000000000b00842300000000000000000000000000000000000000000b00663c00000000000000000000000000000000000000000b00ad3f00000000000000000000000000000000000000000b008f3600000000000000000000000000000000000000000b00f60000000000000000000000000000000000000000000b003a0800000000000000000000000000000000000000000b00ba0e00000000000000000000000000000000000000000b00801000000000000000000000000000000000000000000b00861000000000000000000000000000000000000000000b005a2700000000000000000000000000000000000000000b009b3900000000000000000000000000000000000000000b00b50c00000000000000000000000000000000000000000b00804000000000000000000000000000000000000000000b00901000000000000000000000000000000000000000000b00b84600000000000000000000000000000000000000000b00712e00000000000000000000000000000000000000000b00752e00000000000000000000000000000000000000000b00ff1c00000000000000000000000000000000000000000b00304a00000000000000000000000000000000000000000b005e4300000000000000000000000000000000000000000b001c1f00000000000000000000000000000000000000000b00294a00000000000000000000000000000000000000000b00790700000000000000000000000000000000000000000b00781200000000000000000000000000000000000000000b000c0000000000000000000000000000000000000000000b005f4500000000000000000000000000000000000000000b00441600000000000000000000000000000000000000000b00590000000000000000000000000000000000000000000b00ef1a00000000000000000000000000000000000000000b00fe0500000000000000000000000000000000000000000b00db2500000000000000000000000000000000000000000b00461300000000000000000000000000000000000000000b002c2200000000000000000000000000000000000000000b002d0800000000000000000000000000000000000000000b00934500000000000000000000000000000000000000000b00ca2000000000000000000000000000000000000000000b00cc4600000000000000000000000000000000000000000b00db2000000000000000000000000000000000000000000b00080000000000000000000000000000000000000000000b00760a00000000000000000000000000000000000000000b00e51900000000000000000000000000000000000000000b00270e00000000000000000000000000000000000000000b00524300000000000000000000000000000000000000000b00be1e00000000000000000000000000000000000000000b00790800000000000000000000000000000000000000000b00441900000000000000000000000000000000000000000b00d03d00000000000000000000000000000000000000000b00fd1200000000000000000000000000000000000000000b00242a00000000000000000000000000000000000000000b00d20100000000000000000000000000000000000000000b00a04800000000000000000000000000000000000000000b00394a00000000000000000000000000000000000000000b001f0100000000000000000000000000000000000000000b00331a00000000000000000000000000000000000000000b00cf2f00000000000000000000000000000000000000000b00702600000000000000000000000000000000000000000b00b00b00000000000000000000000000000000000000000b000b4200000000000000000000000000000000000000000b00e22b00000000000000000000000000000000000000000b00dd2f00000000000000000000000000000000000000000b00b60a00000000000000000000000000000000000000000b006b3d00000000000000000000000000000000000000000b00a53c00000000000000000000000000000000000000000b00b92900000000000000000000000000000000000000000b00d63600000000000000000000000000000000000000000b00dc0e00000000000000000000000000000000000000000b00f82900000000000000000000000000000000000000000b00702100000000000000000000000000000000000000000b00b22100000000000000000000000000000000000000000b00513600000000000000000000000000000000000000000b00f73300000000000000000000000000000000000000000b00b02700000000000000000000000000000000000000000b00d54600000000000000000000000000000000000000000b00f60c00000000000000000000000000000000000000000b00082a00000000000000000000000000000000000000000b00fd3300000000000000000000000000000000000000000b00393400000000000000000000000000000000000000000b000a0400000000000000000000000000000000000000000b00473d00000000000000000000000000000000000000000b00bb3000000000000000000000000000000000000000000b00240100000000000000000000000000000000000000000b00460500000000000000000000000000000000000000000b005f4700000000000000000000000000000000000000000b002d4b00000000000000000000000000000000000000000b00674700000000000000000000000000000000000000000b00be2600000000000000000000000000000000000000000b00642c00000000000000000000000000000000000000000b003a3200000000000000000000000000000000000000000b00684500000000000000000000000000000000000000000b00673a00000000000000000000000000000000000000000b00101a00000000000000000000000000000000000000000b00b73100000000000000000000000000000000000000000b005b0e00000000000000000000000000000000000000000b007c2b00000000000000000000000000000000000000000b00441400000000000000000000000000000000000000000b006e4400000000000000000000000000000000000000000b00034700000000000000000000000000000000000000000b00f00c00000000000000000000000000000000000000000b00ec0000000000000000000000000000000000000000000b00df1800000000000000000000000000000000000000000b00f43300000000000000000000000000000000000000000b00e32200000000000000000000000000000000000000000b00d43800000000000000000000000000000000000000000b002e2900000000000000000000000000000000000000000b00464400000000000000000000000000000000000000000b000a2f00000000000000000000000000000000000000000b007f3700000000000000000000000000000000000000000b00624900000000000000000000000000000000000000000b00192a00000000000000000000000000000000000000000b00cc0800000000000000000000000000000000000000000b00330800000000000000000000000000000000000000000b00b43000000000000000000000000000000000000000000b007d0e00000000000000000000000000000000000000000b00370500000000000000000000000000000000000000000b00b44300000000000000000000000000000000000000000b00903a00000000000000000000000000000000000000000b00ba0300000000000000000000000000000000000000000b00334100000000000000000000000000000000000000000b00910600000000000000000000000000000000000000000b00f50d00000000000000000000000000000000000000000b002c3f00000000000000000000000000000000000000000b006c3900000000000000000000000000000000000000000b00662d00000000000000000000000000000000000000000b00f64600000000000000000000000000000000000000000b00664600000000000000000000000000000000000000000b008c4b00000000000000000000000000000000000000000b00e62800000000000000000000000000000000000000000b00cc1500000000000000000000000000000000000000000b00fd2d00000000000000000000000000000000000000000b00113d00000000000000000000000000000000000000000b00e31100000000000000000000000000000000000000000b00450f00000000000000000000000000000000000000000b005f3100000000000000000000000000000000000000000b00243000000000000000000000000000000000000000000b00154200000000000000000000000000000000000000000b00a41900000000000000000000000000000000000000000b00152600000000000000000000000000000000000000000b00fc4400000000000000000000000000000000000000000b00303200000000000000000000000000000000000000000b00c20200000000000000000000000000000000000000000b00d41300000000000000000000000000000000000000000b00ec0400000000000000000000000000000000000000000b00f71100000000000000000000000000000000000000000b00ae4700000000000000000000000000000000000000000b00453200000000000000000000000000000000000000000b00801800000000000000000000000000000000000000000b00cd0600000000000000000000000000000000000000000b00eb3b00000000000000000000000000000000000000000b001a3000000000000000000000000000000000000000000b00bc3e00000000000000000000000000000000000000000b005b0900000000000000000000000000000000000000000b006a2600000000000000000000000000000000000000000b00c01700000000000000000000000000000000000000000b00632200000000000000000000000000000000000000000b00892b00000000000000000000000000000000000000000b00071000000000000000000000000000000000000000000a00f00c00000000000000000000000000000000000000000a00200d00000000000000000000000000000000000000000a00500d00000000000000000000000000000000000000000b008c0600000000000000000000000000000000000000000b00173500000000000000000000000000000000000000000b00db2c00000000000000000000000000000000000000000b00091800000000000000000000000000000000000000000b00121800000000000000000000000000000000000000000b000e2d00000000000000000000000000000000000000000b004c1500000000000000000000000000000000000000000b00b94400000000000000000000000000000000000000000300a84201000000000000000000000000000000000000000300b642010000000000000000000000000000000000000003007877010000000000000000000000000000000000000003007a7701000000000000000000000000000000000000000300bc7801000000000000000000000000000000000000000300a07a01000000000000000000000000000000000000000300f67a010000000000000000000000000000000000000003006e7e010000000000000000000000000000000000000003007c7e01000000000000000000000000000000000000000300fa7f010000000000000000000000000000000000000003000c80010000000000000000000000000000000000000003001e80010000000000000000000000000000000000000003002c80010000000000000000000000000000000000000003003a8001000000000000000000000000000000000000000300488001000000000000000000000000000000000000000300b880010000000000000000000000000000000000000003007482010000000000000000000000000000000000000003002883010000000000000000000000000000000000000003006083010000000000000000000000000000000000000003006a83010000000000000000000000000000000000000003002084010000000000000000000000000000000000000003005a84010000000000000000000000000000000000000003007a8501000000000000000000000000000000000000000300128601000000000000000000000000000000000000000300208601000000000000000000000000000000000000000300368601000000000000000000000000000000000000000300d8860100000000000000000000000000000000000000030048870100000000000000000000000000973800000400f1ff000000000000000000000000000000009d38000000000300eea40100000000000000000000000000a038000000000300bca50100000000000000000000000000a338000000000300e4a90100000000000000000000000000a6380000000003000aaa0100000000000000000000000000a938000000000300baa50100000000000000000000000000ad38000000000300aaa50100000000000000000000000000b138000000000300e0a90100000000000000000000000000b63800000000030098a60100000000000000000000000000bb38000000000300e0a50100000000000000000000000000c03800000000030082a80100000000000000000000000000c538000000000300dca50100000000000000000000000000ca38000000000300aca60100000000000000000000000000cf3800000000030058a60100000000000000000000000000d43800000000030016a60100000000000000000000000000d9380000000003001aa90100000000000000000000000000de3800000000030026a60100000000000000000000000000e3380000000003007ea60100000000000000000000000000e8380000000003008aa60100000000000000000000000000ed380000000003006ca80100000000000000000000000000f23800000000030060a70100000000000000000000000000f7380000000003004aa90100000000000000000000000000fc380000000003008ca801000000000000000000000000000139000000000300f6a601000000000000000000000000000639000000000300faa701000000000000000000000000000b3900000000030042a80100000000000000000000000000103900000000030068a8010000000000000000000000000015390000000003008ea601000000000000000000000000001a39000000000300aea801000000000000000000000000001f3900000000030024a90100000000000000000000000000243900000000030074a901000000000000000000000000002939000000000300f4a501000000000000000000000000002e39000000000300faa901000000000000000000000000003439000000000300fea901000000000000000000000000003a39000000000300e6a901000000000000000000000000004039000000000300eaaa01000000000000000000000000004639000000000300caab01000000000000000000000000004c39000000000300eeaa0100000000000000000000000000523900000000030056ab01000000000000000000000000005839000000000300d0ab01000000000000000000000000005e39000000000300ccab010000000000000000000000000064390000000003006caa01000000000000000000000000006a3900000000030040ab01000000000000000000000000007039000000000300e6ab010000000000000000000000000076390000000003000cab01000000000000000000000000007c3900000000030006ab01000000000000000000000000008239000000000300d6ab010000000000000000000000000088390000000003002aab01000000000000000000000000008e39000000000300eaab010000000000000000000000000094390000000003006eab01000000000000000000000000009a3900000000030068ab0100000000000000000000000000a039000000000300daab0100000000000000000000000000a63900000000030096ab0100000000000000000000000000ac39000000000300b8ab0100000000000000000000000000b239000000000300b6ab0100000000000000000000000000b839000000000300b2ab0100000000000000000000000000be3900000000030020ab0100000000000000000000000000c43900000000030080ab0100000000000000000000000000e039000002020300eea4010000000000ce00000000000000e739000002020300bca50100000000002804000000000000ee39000002020300e4a90100000000002600000000000000f5390000020203000aaa010000000000e601000000000000ca39000012000300ea26010000000000181b000000000000d939000010000300d4260100000000000000000000000000002e726f64617461002e65685f6672616d65002e74657874002e7364617461002e64617461002e627373002e64656275675f616262726576002e64656275675f696e666f002e64656275675f6172616e676573002e64656275675f72616e676573002e64656275675f737472002e64656275675f7075626e616d6573002e64656275675f7075627479706573002e72697363762e61747472696275746573002e64656275675f6c696e65002e636f6d6d656e74002e73796d746162002e7368737472746162002e73747274616200007374616b652e643261633065616565393339383164632d6367752e30002e4c706372656c5f686930005f5a4e37636b625f73746433656e7634415247563137683036373561626564353032343439613545005f5a4e35616c6c6f63377261775f7665633139526177566563244c54245424432441244754243131616c6c6f636174655f696e3137683961373435623837316432623838663945002e4c706372656c5f686931002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e343330002e4c706372656c5f686933002e4c706372656c5f686932005f5a4e34636f726533707472353564726f705f696e5f706c616365244c54246d6f6c6563756c652e2e6572726f722e2e566572696669636174696f6e4572726f72244754243137683936383830623737653965663033383845005f5f727573745f6465616c6c6f63005f5a4e39305f244c54247574696c2e2e6572726f722e2e4572726f72247532302461732475323024636f72652e2e636f6e766572742e2e46726f6d244c5424636b625f7374642e2e6572726f722e2e5379734572726f7224475424244754243466726f6d3137686233643163343538633564356263343545002e4c706372656c5f686934002e4c706372656c5f686935002e4c706372656c5f686936005f5a4e34636f726535736c69636535696e64657837345f244c5424696d706c2475323024636f72652e2e6f70732e2e696e6465782e2e496e646578244c542449244754242475323024666f72247532302424753562245424753564242447542435696e6465783137683064326565363561653136626361336545005f5a4e3131315f244c5424616c6c6f632e2e7665632e2e566563244c54245424475424247532302461732475323024616c6c6f632e2e7665632e2e737065635f66726f6d5f697465725f6e65737465642e2e5370656346726f6d497465724e6573746564244c5424542443244924475424244754243966726f6d5f697465723137683032353562336632346332623633633445005f5a4e35616c6c6f63337665633136566563244c542454244324412447542434707573683137683832346530366138613965323339383745005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f7233616e793137683031323866356465313834336464653445002e4c706372656c5f686938002e4c706372656c5f686937005f5a4e3130325f244c5424636b625f7374616e64616c6f6e655f74797065732e2e67656e6572617465642e2e626c6f636b636861696e2e2e42797465735265616465722475323024617324753230246d6f6c6563756c652e2e7072656c7564652e2e52656164657224475424367665726966793137683135663233383466353032373265326345005f5a4e386d6f6c6563756c6535627974657335427974657335736c6963653137683339643866386561613338343133646245002e4c706372656c5f686939002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e3936002e4c706372656c5f68693130002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e3234005f5a4e386d6f6c6563756c6535627974657335427974657335736c6963653137683133633337653065643765643238336345005f5a4e39385f244c54246d6f6c6563756c65322e2e7265616465722e2e437572736f72247532302461732475323024636f72652e2e636f6e766572742e2e46726f6d244c5424616c6c6f632e2e7665632e2e566563244c542475382447542424475424244754243466726f6d3137686365383937663564613837343036643045005f5a4e396d6f6c6563756c65323672656164657236437572736f723135736c6963655f62795f6f66667365743137683635646335653064333235363034343945005f5a4e396d6f6c6563756c6532367265616465723130385f244c5424696d706c2475323024636f72652e2e636f6e766572742e2e46726f6d244c54246d6f6c6563756c65322e2e7265616465722e2e437572736f72244754242475323024666f722475323024616c6c6f632e2e7665632e2e566563244c5424753824475424244754243466726f6d3137683965653331373661666261663535343545005f5a4e36345f244c5424616c6c6f632e2e72632e2e5263244c54245424475424247532302461732475323024636f72652e2e6f70732e2e64726f702e2e44726f70244754243464726f703137683663346239333364656266363135663545002e4c706372656c5f68693136002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e383436002e4c706372656c5f68693138002e4c706372656c5f68693137002e4c706372656c5f68693139002e4c706372656c5f68693230002e4c706372656c5f68693231002e4c706372656c5f68693233002e4c706372656c5f68693232005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243135636f70795f66726f6d5f736c69636531376c656e5f6d69736d617463685f6661696c3137686531663934356265353831313135613845002e4c706372656c5f68693131007374722e342e3436005f5a4e34636f72653970616e69636b696e673570616e69633137686437373538656430613265383739363145005f5a4e39385f244c5424636b625f7374642e2e686967685f6c6576656c2e2e517565727949746572244c54244624475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137686231366136333531633137303061613745005f5a4e37636b625f7374643130686967685f6c6576656c31346c6f61645f63656c6c5f646174613137686438663961623933373437336639633645005f5a4e396d6f6c6563756c65323672656164657236437572736f7232307461626c655f736c6963655f62795f696e6465783137686232343839353738643638326165663045005f5a4e347574696c3668656c70657231356765745f7363726970745f686173683137683861333134336361336163636135633445005f5a4e37636b625f7374643130686967685f6c6576656c31396c6f61645f63656c6c5f6c6f636b5f686173683137686238376330343133623735373432633545005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f72656164657237547970654964733134787564745f747970655f686173683137686334653636633566343738343237356145005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f726561646572375479706549647331397374616b655f736d745f636f64655f686173683137683939313230643232643561376161363745005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f726561646572375479706549647331377374616b655f736d745f747970655f69643137683133613730383736373561386135323245005f5a4e347574696c3668656c70657232376765745f63656c6c5f636f756e745f62795f747970655f686173683137683636366663636666636434353161366445005f5a4e347574696c3668656c7065723230636865636b5f787564745f747970655f686173683137683036636334386162663931333435343345005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231355374616b65417443656c6c4461746131366d657461646174615f747970655f69643137683136353731366261626264366365656645005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f72656164657237547970654964733138636865636b706f696e745f747970655f69643137683062376537323033303666383865346345005f5a4e347574696c3668656c70657232316765745f787564745f62795f747970655f686173683137686133323939383965653034636166616145002e4c706372656c5f68693238007374722e302e333235002e4c706372656c5f68693132002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3436002e4c706372656c5f68693133002e4c616e6f6e2e65383134633736363361666663333138633766356639363865643531663662352e3139002e4c706372656c5f68693134002e4c706372656c5f68693135005f5a4e34636f726536726573756c743133756e777261705f6661696c65643137683030653934303161326339653536633045005f5a4e347574696c3668656c70657233306765745f7374616b655f61745f646174615f62795f6c6f636b5f686173683137683536356232313136353933333665623945005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231345374616b65496e666f44656c7461313169735f696e6372656173653137683166386136356661303836623163316645005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231355374616b65417443656c6c446174613564656c74613137683762333332613765343438316530613845005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231345374616b65496e666f44656c746136616d6f756e743137683736303137613463316430633135626445005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231345374616b65496e666f44656c74613138696e61756775726174696f6e5f65706f63683137683538323561303933383837366165313345005f5a4e347574696c3668656c70657231376765745f63757272656e745f65706f63683137683433313039626562306665666534313945002e4c706372656c5f68693236002e4c706372656c5f68693237002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3438002e4c706372656c5f68693234002e4c706372656c5f68693235002e4c616e6f6e2e36633237623166666234666234346562313164656530663863336331326232322e32002e4c706372656c5f68693239002e4c706372656c5f68693330002e4c706372656c5f68693331002e4c706372656c5f68693332002e4c706372656c5f68693333002e4c706372656c5f68693334002e4c706372656c5f68693335002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e34002e4c706372656c5f68693336007374722e30002e4c706372656c5f68693337007374722e31002e4c706372656c5f68693430002e4c706372656c5f68693339002e4c706372656c5f6869333800727573745f626567696e5f756e77696e64005f5a4e37636b625f7374643873797363616c6c73366e617469766534657869743137683163616638653234666532613530323145005f5f72675f616c6c6f63005f5a4e3130365f244c542462756464795f616c6c6f632e2e6e6f6e5f746872656164736166655f616c6c6f632e2e4e6f6e54687265616473616665416c6c6f63247532302461732475323024636f72652e2e616c6c6f632e2e676c6f62616c2e2e476c6f62616c416c6c6f632447542435616c6c6f633137683966656332343337626566343266383945005f5f72675f6465616c6c6f63005f5a4e3130365f244c542462756464795f616c6c6f632e2e6e6f6e5f746872656164736166655f616c6c6f632e2e4e6f6e54687265616473616665416c6c6f63247532302461732475323024636f72652e2e616c6c6f632e2e676c6f62616c2e2e476c6f62616c416c6c6f6324475424376465616c6c6f633137686530336235656339643238613732396445005f5f72675f7265616c6c6f63005f5f72675f616c6c6f635f7a65726f6564005f5a4e35616c6c6f63377261775f766563313763617061636974795f6f766572666c6f773137683736396433373734353939336431626545005f5a4e34636f72653970616e69636b696e67313870616e69635f6e6f756e77696e645f666d743137683133386130386530383963323036303445005f5f72646c5f6f6f6d002e4c706372656c5f68693431002e4c706372656c5f68693432002e4c706372656c5f68693433002e4c706372656c5f68693434002e4c706372656c5f68693435002e4c706372656c5f68693436002e4c706372656c5f68693437002e4c706372656c5f68693438005f5a4e396d6f6c6563756c65323672656164657238355f244c5424696d706c2475323024636f72652e2e636f6e766572742e2e46726f6d244c54246d6f6c6563756c65322e2e7265616465722e2e437572736f72244754242475323024666f7224753230247538244754243466726f6d3137686461653235633931336631613435396545002e4c706372656c5f68693439002e4c706372656c5f68693530002e4c706372656c5f68693531002e4c706372656c5f68693532005f5a4e396d6f6c6563756c65323672656164657238365f244c5424696d706c2475323024636f72652e2e636f6e766572742e2e46726f6d244c54246d6f6c6563756c65322e2e7265616465722e2e437572736f72244754242475323024666f722475323024753634244754243466726f6d3137686232663035653938653831303635333145002e4c706372656c5f68693533002e4c706372656c5f68693534002e4c706372656c5f68693535002e4c706372656c5f68693536002e4c706372656c5f68693537002e4c706372656c5f68693538005f5a4e3131626c616b6532625f7265663131626c616b6532625f7265663138626c616b6532625f696e69745f706172616d3137683431613831343963666239633164343445002e4c706372656c5f68693539005f5a4e3131626c616b6532625f7265663131626c616b6532625f7265663130626c616b6532625f49563137686532356438333932346363316638393145005f5a4e3131626c616b6532625f7265663131626c616b6532625f7265663134626c616b6532625f7570646174653137683337646637643338333264666265336545005f5a4e3131626c616b6532625f7265663131626c616b6532625f7265663136626c616b6532625f636f6d70726573733137683531363361326435303733336262323945002e4c43504931395f30002e4c43504931395f31002e4c43504931395f32002e4c43504931395f33002e4c43504931395f34002e4c43504931395f35002e4c43504931395f36002e4c43504931395f37002e4c706372656c5f68693630002e4c706372656c5f68693631002e4c706372656c5f68693632002e4c706372656c5f68693633002e4c706372656c5f68693634002e4c706372656c5f68693635002e4c706372656c5f68693636002e4c706372656c5f68693637005f5a4e313162756464795f616c6c6f63313162756464795f616c6c6f6331304275646479416c6c6f63336e65773137683039343964346234353436656265666245005f5a4e313162756464795f616c6c6f63313162756464795f616c6c6f6337726f756e6475703137686533656266373734346663663366363345002e4c706372656c5f68693735007374722e342e3336005f5a4e313162756464795f616c6c6f63313162756464795f616c6c6f63366e626c6f636b3137683537623963376462363561386133343745005f5a4e313162756464795f616c6c6f63313162756464795f616c6c6f6331304275646479416c6c6f633131626c6f636b5f696e6465783137683333633165376336333564613363643945005f5a4e34636f7265366f7074696f6e31336578706563745f6661696c65643137686332333330616533386638616564396545002e4c706372656c5f68693830002e4c706372656c5f68693736002e4c706372656c5f68693737002e4c706372656c5f68693638002e4c706372656c5f68693730007374722e322e3337002e4c706372656c5f68693731007374722e332e3338002e4c706372656c5f68693732002e4c706372656c5f68693733007374722e312e3335002e4c706372656c5f68693734002e4c706372656c5f68693831002e4c706372656c5f68693738007374722e302e3334002e4c706372656c5f68693639002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3135002e4c706372656c5f68693832002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3238005f5a4e34636f72653970616e69636b696e67313370616e69635f646973706c61793137683538303536323433613031393534316645002e4c706372656c5f68693739002e4c706372656c5f68693833002e4c706372656c5f68693834002e4c706372656c5f68693835002e4c706372656c5f68693836002e4c706372656c5f68693837002e4c706372656c5f68693839002e4c706372656c5f68693930002e4c706372656c5f68693838002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3338005f5a4e313162756464795f616c6c6f633130666173745f616c6c6f633946617374416c6c6f63336e65773137683239303962396561363461333531383845002e4c706372656c5f68693932002e4c706372656c5f68693931002e4c706372656c5f68693933002e4c706372656c5f68693934005f5a4e357374616b6535414c4c4f433137683735313734646435353830643734633445002e4c706372656c5f68693938002e4c706372656c5f6869313033002e4c706372656c5f6869313034002e4c706372656c5f6869313031002e4c706372656c5f6869313035002e4c706372656c5f6869313036002e4c706372656c5f6869313032002e4c706372656c5f68693937002e4c706372656c5f68693939002e4c706372656c5f6869313030002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e32002e4c706372656c5f68693935002e4c706372656c5f68693936002e4c706372656c5f6869313037002e4c706372656c5f6869313038002e4c706372656c5f6869313039002e4c706372656c5f6869313133002e4c706372656c5f6869313132002e4c706372656c5f6869313136002e4c706372656c5f6869313138002e4c706372656c5f6869313139002e4c706372656c5f6869313230002e4c706372656c5f6869313137002e4c706372656c5f6869313130002e4c706372656c5f6869313131002e4c706372656c5f6869313134002e4c706372656c5f6869313135005f5a4e35616c6c6f63377261775f7665633139526177566563244c54245424432441244754243131616c6c6f636174655f696e3137683334393639363464643031633234363645005f5a4e35616c6c6f63377261775f7665633139526177566563244c542454244324412447542437726573657276653231646f5f726573657276655f616e645f68616e646c653137686234636364626536643135363830353445002e4c706372656c5f6869313231007374722e302e3434005f5f727573745f616c6c6f63005f5f727573745f616c6c6f635f6572726f725f68616e646c6572005f5a4e35616c6c6f63377261775f7665633139526177566563244c5424542443244124475424313467726f775f616d6f7274697a65643137683131313435313531653037646531613245005f5a4e35616c6c6f63377261775f766563313166696e6973685f67726f773137683362363537323731663362336132663345005f5a4e35616c6c6f63377261775f7665633139526177566563244c54245424432441244754243136726573657276655f666f725f707573683137683364383734353931323332303230376445002e4c706372656c5f6869313232002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e313734002e4c706372656c5f6869313233002e4c706372656c5f6869313234005f5a4e36315f244c5424636b625f7374642e2e6572726f722e2e5379734572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683863383033303266623836336136303845002e4c706372656c5f6869313235002e4c4a544933395f30002e4c424233395f31002e4c706372656c5f6869313236002e4c616e6f6e2e34313466363731613135666237623063306532636261396133343630323939342e3339002e4c424233395f32002e4c706372656c5f6869313237002e4c616e6f6e2e34313466363731613135666237623063306532636261396133343630323939342e3338002e4c424233395f33002e4c706372656c5f6869313238002e4c616e6f6e2e34313466363731613135666237623063306532636261396133343630323939342e3336002e4c706372656c5f6869313239002e4c616e6f6e2e34313466363731613135666237623063306532636261396133343630323939342e3337002e4c424233395f34002e4c706372656c5f6869313330002e4c424233395f36002e4c706372656c5f6869313331002e4c616e6f6e2e34313466363731613135666237623063306532636261396133343630323939342e3333002e4c706372656c5f6869313332002e4c616e6f6e2e34313466363731613135666237623063306532636261396133343630323939342e3334005f5a4e34636f726533666d7439466f726d6174746572323564656275675f7475706c655f6669656c64315f66696e6973683137683963326264643732306464613133376545005f5a4e34636f726533707472323864726f705f696e5f706c616365244c542424524624753634244754243137683536663832373834643464373061633345005f5a4e37636b625f7374643130686967685f6c6576656c31396c6f61645f63656c6c5f747970655f686173683137686661353738353337303831333261613945005f5a4e34636f7265336f70733866756e6374696f6e36466e4f6e63653963616c6c5f6f6e63653137683331326365396462383432326365623645005f5a4e34636f72653370747231303264726f705f696e5f706c616365244c542424524624636f72652e2e697465722e2e61646170746572732e2e636f706965642e2e436f70696564244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c542475382447542424475424244754243137683465633534623435323134663763393045002e4c43504934385f30005f5a4e34636f726533666d74336e756d33696d7037666d745f7536343137683238366534643532373433386334363745002e4c706372656c5f6869313333002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333234002e4c706372656c5f6869313334002e4c706372656c5f6869313335002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3233005f5a4e34636f726533666d7439466f726d617474657231327061645f696e74656772616c3137686238656639343965396131613633346545005f5a4e34636f726533666d7439466f726d617474657231327061645f696e74656772616c313277726974655f7072656669783137683834663538656430383761336264393345002e4c43504935315f30002e4c43504935315f31005f5a4e34636f726533666d7439466f726d6174746572337061643137683433336537613934646232626438653245002e4c706372656c5f6869313336002e4c706372656c5f6869313337005f5a4e34636f726533666d743577726974653137683537653362636463656237646630393145002e4c706372656c5f6869313338005f5a4e36305f244c5424636f72652e2e63656c6c2e2e426f72726f774572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137686163386261333334363731373261333845002e4c706372656c5f6869313339002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e313730005f5a4e36335f244c5424636f72652e2e63656c6c2e2e426f72726f774d75744572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683636336332373865383138373636393045002e4c706372656c5f6869313430002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e313731005f5a4e34636f726533666d74336e756d35335f244c5424696d706c2475323024636f72652e2e666d742e2e4c6f7765724865782475323024666f7224753230246936342447542433666d743137686632356530653835343735353364373145002e4c706372656c5f6869313431002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333232002e4c43504936305f30002e4c43504936305f31002e4c43504936305f32005f5a4e36385f244c5424636f72652e2e666d742e2e6275696c646572732e2e50616441646170746572247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f7374723137686539366438303337316562386433343445002e4c706372656c5f6869313432002e4c706372656c5f6869313433002e4c706372656c5f6869313434002e4c706372656c5f6869313435005f5a4e34636f726533666d74355772697465313077726974655f636861723137686664666234386663643336373461323845005f5a4e34636f726533666d743557726974653977726974655f666d743137683364623431343565346436363932376245002e4c706372656c5f6869313436002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333237005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f7374723137683865303931326361326264646233386345005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e577269746524475424313077726974655f636861723137683239666437616639333939643762333645005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f666d743137683565373464633863623261616161323645002e4c706372656c5f6869313437005f5a4e34636f726533666d74386275696c64657273313044656275675475706c65356669656c643137686134393061356537663734366534656245002e4c706372656c5f6869313439002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e323933002e4c706372656c5f6869313530002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333030002e4c706372656c5f6869313438002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333031002e4c706372656c5f6869313531002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e323839002e4c706372656c5f6869313532002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e323932002e4c706372656c5f6869313534002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333032002e4c706372656c5f6869313533002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e313537005f5a4e34325f244c54242452462454247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137686332303631326561373836393861653445002e4c706372656c5f6869313535002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333337005f5a4e36375f244c5424636f72652e2e61727261792e2e54727946726f6d536c6963654572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683532646436363362353834636335356645002e4c706372656c5f6869313536002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e353537002e4c706372656c5f6869313537002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e353333002e4c706372656c5f6869313539002e4c706372656c5f6869313538005f5a4e34636f726533666d74336e756d35335f244c5424696d706c2475323024636f72652e2e666d742e2e55707065724865782475323024666f7224753230246936342447542433666d743137683464336136353331313038303933376445002e4c706372656c5f6869313630005f5a4e3133325f244c5424616c6c6f632e2e7665632e2e566563244c5424542443244124475424247532302461732475323024616c6c6f632e2e7665632e2e737065635f657874656e642e2e53706563457874656e64244c54242452462454244324636f72652e2e736c6963652e2e697465722e2e49746572244c5424542447542424475424244754243131737065635f657874656e643137683464663561353366366631653763336445005f5a4e35616c6c6f63377261775f7665633139526177566563244c542454244324412447542437726573657276653231646f5f726573657276655f616e645f68616e646c653137686332663335393562613638613033633645005f5f727573745f7265616c6c6f63005f5a4e34325f244c54242452462454247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683431323134373832613466363464656645005f5f727573745f616c6c6f635f7a65726f6564005f5a4e35616c6c6f63337665633136566563244c54245424432441244754243131657874656e645f776974683137683935323361376565386561616133316645005f5a4e35616c6c6f63377261775f7665633139526177566563244c542454244324412447542437726573657276653231646f5f726573657276655f616e645f68616e646c653137686534386235666233366361343936633545005f5a4e35616c6c6f63377261775f766563313166696e6973685f67726f773137686465323762646133633136313431313345005f5a4e396d6f6c6563756c65323672656164657237726561645f61743137686436323832346538376630396538383045002e4c706372656c5f6869313730007374722e312e323830002e4c706372656c5f6869313633002e4c706372656c5f6869313634002e4c706372656c5f6869313631002e4c706372656c5f6869313632002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e31002e4c706372656c5f6869313639002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3136002e4c706372656c5f6869313731002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3139002e4c706372656c5f6869313635002e4c706372656c5f6869313636002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e36002e4c706372656c5f6869313637002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3132002e4c706372656c5f6869313638002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3134005f5a4e36315f244c54246d6f6c6563756c65322e2e7265616465722e2e4572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683238346238363235356264316239336545002e4c706372656c5f6869313732002e4c7377697463682e7461626c652e5f5a4e36315f244c54246d6f6c6563756c65322e2e7265616465722e2e4572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683238346238363235356264316239336545002e4c706372656c5f6869313733002e4c7377697463682e7461626c652e5f5a4e36315f244c54246d6f6c6563756c65322e2e7265616465722e2e4572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d7431376832383462383632353562643162393365452e333731005f5a4e396d6f6c6563756c65323672656164657236437572736f723876616c69646174653137683930306131623931383065653939313845002e4c706372656c5f6869313736002e4c706372656c5f6869313734002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e32002e4c706372656c5f6869313735002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e33002e4c706372656c5f6869313737002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3238005f5a4e396d6f6c6563756c65323672656164657236437572736f723133756e7061636b5f6e756d6265723137683635326430373132666263326536343145002e4c706372656c5f6869313738002e4c706372656c5f6869313739002e4c706372656c5f6869313830002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3331002e4c706372656c5f6869313831002e4c706372656c5f6869313839002e4c706372656c5f6869313832002e4c706372656c5f6869313833002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3335002e4c706372656c5f6869313834002e4c706372656c5f6869313838002e4c706372656c5f6869313835002e4c706372656c5f6869313836002e4c706372656c5f6869313837002e4c706372656c5f6869313930002e4c706372656c5f6869313931002e4c706372656c5f6869313932002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3430002e4c706372656c5f6869313933002e4c706372656c5f6869313934002e4c706372656c5f6869313935002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3538002e4c706372656c5f6869313936002e4c706372656c5f6869313937002e4c706372656c5f6869313938002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3634005f5a4e36395f244c5424616c6c6f632e2e7665632e2e566563244c54247538244754242475323024617324753230246d6f6c6563756c65322e2e7265616465722e2e526561642447542434726561643137683538323363346134366134643066373445002e4c706372656c5f6869313939002e4c706372656c5f6869323030002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3638005f5a4e34636f726533707472343664726f705f696e5f706c616365244c5424616c6c6f632e2e7665632e2e566563244c5424753824475424244754243137683139303635656264313265376238616645002e4c706372656c5f6869323031005f5a4e3130325f244c5424636f72652e2e697465722e2e61646170746572732e2e6d61702e2e4d6170244c5424492443244624475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424387472795f666f6c643137686134643535656336343238393364643045002e4c706372656c5f6869323035002e4c706372656c5f6869323034002e4c706372656c5f6869323032002e4c706372656c5f6869323033002e4c706372656c5f6869323036002e4c4a54493130305f30002e4c42423130305f31002e4c42423130305f32002e4c42423130305f33002e4c42423130305f34002e4c42423130305f35002e4c706372656c5f6869323134002e4c706372656c5f6869323039007374722e322e3433002e4c706372656c5f6869323130002e4c706372656c5f6869323131002e4c706372656c5f6869323132002e4c706372656c5f6869323133002e4c706372656c5f6869323037002e4c706372656c5f6869323038002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3437002e4c706372656c5f6869323136002e4c706372656c5f6869323135002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e313134002e4c706372656c5f6869323137002e4c706372656c5f6869323138002e4c706372656c5f6869323139002e4c706372656c5f6869323230002e4c706372656c5f6869323231002e4c706372656c5f6869323232002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e313139002e4c706372656c5f6869323233005f5a4e357374616b6531315f42554444595f484541503137683862313032653565633363313635316445005f5a4e357374616b6531375f46495845445f424c4f434b5f484541503137686132366633373037356664663339316245002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3134002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3237002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3732002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3733002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3734002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3735002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3736002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3737002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3738002e4c6c696e655f7461626c655f737461727430002e4c6c696e655f7461626c655f737461727431006c69622e63002478002478002478002478002e4c32002e4c33002e4c3335002e4c3437002e4c3132002e4c3739002e4c3830002e4c3134002e4c3135002e4c3136002e4c3831002e4c3138002e4c3230002e4c3231002e4c3738002e4c3235002e4c3236002e4c3237002e4c3238002e4c3331002e4c3332002e4c3333002e4c3334002e4c3330002e4c3137002e4c3239002e4c3130002e4c313433002e4c313437002e4c313438002e4c313439002e4c323033002e4c313532002e4c323034002e4c313735002e4c313736002e4c313632002e4c323031002e4c313737002e4c313638002e4c313730002e4c313738002e4c313731002e4c313733002e4c313536002e4c313539002e4c313630002e4c313631002e4c313634002e4c323035002e4c313537002e4c313637002e4c313534005f5f636b625f7374645f6d61696e005f7374617274006d656d736574006d656d637079006d656d636d70006d656d6d6f7665000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000120000000000000060010100000000006001000000000000680900000000000000000000000000001000000000000000000000000000000009000000010000000200000000000000c80a010000000000c80a0000000000000c0c00000000000000000000000000000800000000000000000000000000000013000000010000000600000000000000d426010000000000d4160000000000001c8500000000000000000000000000000400000000000000000000000000000019000000010000000300000000000000f0bb010000000000f09b00000000000070000000000000000000000000000000080000000000000000000000000000002000000001000000030000000000000060bc010000000000609c000000000000b8000000000000000000000000000000080000000000000000000000000000002600000008000000030000000000000018bd010000000000189d00000000000000200800000000000000000000000000010000000000000000000000000000002b0000000100000000000000000000000000000000000000189d0000000000002802000000000000000000000000000001000000000000000000000000000000390000000100000000000000000000000000000000000000409f0000000000003f230000000000000000000000000000010000000000000000000000000000004500000001000000000000000000000000000000000000007fc200000000000000020000000000000000000000000000010000000000000000000000000000005400000001000000000000000000000000000000000000007fc40000000000005010000000000000000000000000000001000000000000000000000000000000620000000100000030000000000000000000000000000000cfd40000000000005a4c0000000000000000000000000000010000000000000001000000000000006d00000001000000000000000000000000000000000000002921010000000000481b0000000000000000000000000000010000000000000000000000000000007d0000000100000000000000000000000000000000000000713c01000000000024000000000000000000000000000000010000000000000000000000000000008d0000000300007000000000000000000000000000000000953c0100000000002b000000000000000000000000000000010000000000000000000000000000009f0000000100000000000000000000000000000000000000c03c010000000000791c000000000000000000000000000001000000000000000000000000000000ab000000010000003000000000000000000000000000000039590100000000002300000000000000000000000000000001000000000000000100000000000000b400000002000000000000000000000000000000000000006059010000000000f8e2000000000000130000007309000008000000000000001800000000000000bc0000000300000000000000000000000000000000000000583c020000000000ce00000000000000000000000000000001000000000000000000000000000000c60000000300000000000000000000000000000000000000263d020000000000fd39000000000000000000000000000001000000000000000000000000000000",
      "0x7f454c460201010000000000000000000200f3000100000074360100000000004000000000000000c00f04000000000001000000400038000500400016001400060000000400000040000000000000004000010000000000400001000000000018010000000000001801000000000000080000000000000001000000040000000000000000000000000001000000000000000100000000007426000000000000742600000000000000100000000000000100000005000000742600000000000074360100000000007436010000000000be82010000000000be820100000000000010000000000000010000000600000038a901000000000038c902000000000038c902000000000068010000000000006821080000000000001000000000000051e574640600000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000005ca90100000000006ea901000000000080a901000000000098a9010000000000aea9010000000000383802000000000036380200000000003a380200000000003e38020000000000423802000000000056880200000000000093020000000000009302000000000000930200000000002a8a020000000000009302000000000000930200000000008e8c0200000000004a8e0200000000009a8e020000000000617474656d707420746f206164642077697468206f766572666c6f7700000000ee3601000000000018000000000000000800000000000000c8c6010000000000d8a901000000000000000000000000000100000000000000d0c3010000000000d8a9010000000000010000000000000001000000000000005eca010000000000617474656d707420746f206164642077697468206f766572666c6f770000000008c9bcf367e6096a3ba7ca8485ae67bb2bf894fe72f36e3cf1361d5f3af54fa5d182e6ad7f520e511f6c3e2b8c68059b6bbd41fbabd9831f79217e1319cde05bd8a901000000000000000000000000000100000000000000c2bb010000000000617474656d707420746f207368696674206c6566742077697468206f766572666c6f7700000000000000000000000000617474656d707420746f206d756c7469706c792077697468206f766572666c6f77000000000000000000000000000000617474656d707420746f2073756274726163742077697468206f766572666c6f77000000000000000000000000000000617474656d707420746f2073686966742072696768742077697468206f766572666c6f77000000000000000000000000617474656d707420746f206164642077697468206f766572666c6f776c6561662073697a65206d75737420626520616c69676e20746f20313620627974657300dc0301000000000023000000000000007265717569726573206d6f7265206d656d6f727920737061636520746f20696e697469616c697a65204275646479416c6c6f630000000000100401000000000033000000000000006f7574206f66206d656d6f72790000000000000000000000617474656d707420746f20646976696465206279207a65726f00000000000000617474656d707420746f206164642077697468206f766572666c6f77427974655265616465724279746533325265616465724279746573526561646572000000617474656d707420746f2073756274726163742077697468206f766572666c6f7753637269707452656164657243656c6c496e7075745265616465725769746e65737341726773526561646572556e6b6e6f776e00000000d8a9010000000000080000000000000008000000000000004ac6010000000000456e636f64696e674f766572666c6f7776616c69646174654c656e6774684e6f74456e6f75676800d8a9010000000000080000000000000008000000000000004ac60100000000004974656d4d697373696e67496e6465784f75744f66426f756e64000000000000617474656d707420746f206164642077697468206f766572666c6f7729426f72726f774572726f72426f72726f774d75744572726f725b002eb3010000000000180000000000000008000000000000006ebc0100000000002abe010000000000debe0100000000002020202052656164446174612c0a2c20280a282c0a5d307830303031303230333034303530363037303830393130313131323133313431353136313731383139323032313232323332343235323632373238323933303331333233333334333533363337333833393430343134323433343434353436343734383439353035313532353335343535353635373538353936303631363236333634363536363637363836393730373137323733373437353736373737383739383038313832383338343835383638373838383939303931393239333934393539363937393839392eb30100000000000800000000000000080000000000000016bf01000000000020bf010000000000d6bf01000000000028290000000000002eb301000000000008000000000000000800000000000000bac301000000000054727946726f6d536c6963654572726f72636b622d64656661756c742d68617368616c726561647920626f72726f77656400000000000000d8a901000000000000000000000000000100000000000000c2bb010000000000616c7265616479206d757461626c7920626f72726f776564d8a901000000000000000000000000000100000000000000b0bb010000000000d8a9010000000000010000000000000001000000000000005eca010000000000617474656d707420746f206164642077697468206f766572666c6f77726561645f6174206069662073697a65203c20726561645f6c656e60726561645f6174206069662064732e63616368655f73697a65203e2064732e6d61785f63616368655f73697a6560726561645f617420606966206375722e6f6666736574203c2064732e73746172745f706f696e74207c7c202e2e2e60726561645f61742060696620726561645f706f696e74202b20726561645f6c656e203e2064732e63616368655f73697a656076616c69646174653a2073697a65203e206375722e736f757263652e746f74616c5f73697a65756e7061636b5f6e756d6265726765745f6974656d5f636f756e74636f6e766572745f746f5f753634636f6e766572745f746f5f753136636f6e766572745f746f5f7538636f6e7665727420746f205665633c75383e000000000016d001000000000018000000000000000800000000000000e2ce0100000000004669656c64436f756e744f75744f66426f756e64556e6b6e6f776e4974656d4f6666736574486561646572546f74616c53697a65436f6d6d6f6e617373657274696f6e206661696c65643a20696478203c204341504143495459000000000000000000000000000000000000000000000000000000000000000063616c6c656420604f7074696f6e3a3a756e77726170282960206f6e206120604e6f6e65602076616c7565000000617474656d707420746f206164642077697468206f766572666c6f7700000000617373657274696f6e206661696c65643a206f666673657420213d2030202626206f6666736574203c3d206c656e63616c6c65642060526573756c743a3a756e77726170282960206f6e20616e2060457272602076616c756500000000000000d8a901000000000000000000000000000100000000000000d0c3010000000000d8a90100000000001000000000000000080000000000000046a9010000000000ee3601000000000018000000000000000800000000000000c8c6010000000000617373657274696f6e206661696c65643a20656467652e686569676874203d3d2073656c662e686569676874202d2031617373657274696f6e206661696c65643a2073656c662e686569676874203e2030617373657274696f6e206661696c65643a207372632e6c656e2829203d3d206473742e6c656e2829617373657274696f6e206661696c65643a20656467652e686569676874203d3d2073656c662e6e6f64652e686569676874202d2031617373657274696f6e206661696c65643a20636f756e74203e2030617373657274696f6e206661696c65643a206f6c645f72696768745f6c656e202b20636f756e74203c3d204341504143495459617373657274696f6e206661696c65643a206f6c645f6c6566745f6c656e203e3d20636f756e74696e7465726e616c206572726f723a20656e746572656420756e726561636861626c6520636f6465617373657274696f6e206661696c65643a206f6c645f6c6566745f6c656e202b20636f756e74203c3d204341504143495459617373657274696f6e206661696c65643a206f6c645f72696768745f6c656e203e3d20636f756e74617373657274696f6e206661696c65643a206d6174636820747261636b5f656467655f696478207b5c6e202020204c6566744f7252696768743a3a4c6566742869647829203d3e20696478203c3d206f6c645f6c6566745f6c656e2c5c6e202020204c6566744f7252696768743a3a52696768742869647829203d3e20696478203c3d2072696768745f6c656e2c5c6e7d617373657274696f6e206661696c65643a206e65775f6c6566745f6c656e203c3d204341504143495459617373657274696f6e206661696c65643a20636865636b706f696e745f646174612e69735f6e6f6e652829617373657274696f6e206661696c65643a207374616b655f61745f646174612e69735f6e6f6e652829617373657274696f6e206661696c65643a2077697468647261775f61745f646174612e69735f6e6f6e65282906000000000000000900000000000000060000000000000006000000000000000b000000000000000a000000000000000a000000000000000400000000000000080000000000000004000000000000009c0901000000000093090100000000008d0901000000000087090100000000007c0901000000000072090100000000006809010000000000200601000000000050050100000000001c0601000000000008c9bcf367e6096a2bf894fe72f36e3c1f6c3e2b8c68059b3ba7ca8485ae67bb79217e1319cde05bd182e6ad7f520e51f1361d5f3af54fa56bbd41fbabd9831f1000000000000000017a5200017801011b0c02001c00000018000000be2700006400000000420e2048810188028903920400000010000000380000000228000010000000000000001c0000004c000000fe270000ee00000000420e304a81018802890392049305002c0000006c000000cc280000d404000000420e80035a810188028903920493059406950796089709980a990b9a0c9b0d100000009c000000702d000068000000000e000028000000b0000000c42d0000dc00000000420e6056810188028903920493059406950796089709980a990b0014000000dc000000742e00003000000000420e104281010014000000f40000008c2e00003000000000420e10428101002c0000000c010000a42e00007a01000000420e900158810188028903920493059406950796089709980a990b9a0c00002c0000003c010000ee2f0000aa01000000420ea0015a810188028903920493059406950796089709980a990b9a0c9b0d2c0000006c01000068310000c001000000420ed0015a810188028903920493059406950796089709980a990b9a0c9b0d2c0000009c010000f83200008201000000420eb0015a810188028903920493059406950796089709980a990b9a0c9b0d2c000000cc0100004a3400005002000000420ed0035a810188028903920493059406950796089709980a990b9a0c9b0d2c000000fc0100006a360000c600000000420e6058810188028903920493059406950796089709980a990b9a0c000000300000002c020000003700009025000000440ef00f74810188028903920493059406950796089709980a990b9a0c9b0d420e801210000000600200005c5c00000a000000000e00001000000074020000525c000008000000000000001000000088020000465c000008000000000000001c0000009c0200003a5c00004e00000000420e304a810188028903920493050018000000bc020000685c00003000000000420e20468101880289030010000000d80200007c5c0000080000000000000010000000ec020000705c000008000000000000001000000000030000645c000008000000000000001000000014030000585c0000080000000000000010000000280300004c5c00000a000000000e0000140000003c030000425c00000e00000000420e10428101001400000054030000385c00000e00000000420e1042810100180000006c0300002e5c00005800000000420e40448101880200000018000000880300006a5c00005800000000420e40448101880200000018000000a4030000a65c00005800000000420e40448101880200000018000000c0030000e25c00005800000000420e40448101880200000018000000dc0300001e5d00005800000000420e40448101880200000018000000f80300005a5d00005800000000420e4044810188020000001800000014040000965d00005800000000420e4044810188020000001800000030040000d25d00005800000000420e404481018802000000140000004c0400000e5e00005200000000420e40428101001800000064040000485e00005800000000420e4044810188020000001400000080040000845e00005200000000420e40428101001800000098040000be5e00004e00000000420e30448101880200000018000000b4040000f05e00005800000000420e40448101880200000018000000d00400002c5f00005800000000420e40448101880200000018000000ec040000685f00008600000000420e3046810188028903001800000008050000d25f00004c00000000420e3044810188020000001800000024050000026000004e00000000420e3044810188020000001800000040050000346000009400000000420e604481018802000000180000005c050000ac6000009400000000420e6044810188020000001c0000007805000024610000bc00000000420ee00348810188028903920400001c00000098050000c06100009a00000000420e2048810188028903920400000020000000b80500003a620000dc00000000440e304c8101880289039204930594060000002c000000dc050000f2620000ee1a000000420ef0035a810188028903920493059406950796089709980a990b9a0c9b0d1c0000000c060000b07d0000f000000000420e60488101880289039204000000180000002c060000807e00007c00000000420e9003468101880289032c00000048060000e07e00001404000000420e80015a810188028903920493059406950796089709980a990b9a0c9b0d1000000078060000c48200003c000000000e0000100000008c060000ec8200000a000000000e000010000000a0060000e28200004c000000000e000010000000b40600001a8300004c000000000e000010000000c806000052830000f4000000000e00002c000000dc06000032840000d403000000420eb00158810188028903920493059406950796089709980a990b9a0c00002c0000000c070000d6870000f203000000420ec0015a810188028903920493059406950796089709980a990b9a0c9b0d200000003c070000988b0000d600000000420e504e81018802890392049305940695070018000000600700004a8c00005200000000420e204681018802890300140000007c070000808c00003400000000420e104281010018000000940700009c8c00007400000000420e50468101880289030014000000b0070000f48c00003600000000420e104281010020000000c8070000128d00006c00000000420e304c81018802890392049305940600000010000000ec0700005a8d000022000000000e00001800000000080000688d00003a00000000420e204681018802890300200000001c080000868d0000fc00000000420e404e81018802890392049305940695070010000000400800005e8e000042000000000e000020000000540800008c8e00005000000000420e304c8101880289039204930594060000001c00000078080000b88e00007400000000420e4048810188028903920400000020000000980800000c8f00006400000000420e304c8101880289039204930594060000001c000000bc0800004c8f00008200000000420e2048810188028903920400000028000000dc080000ae8f00009601000000420e900154810188028903920493059406950796089709980a000010000000080900001891000072000000000e0000140000001c090000769100009200000000420e10428101001000000034090000f091000002000000000000001000000048090000de9100003600000000000000240000005c09000000920000c001000000440ee008648101880289039204930594069507960897091800000084090000989300007a00000000420e40448101880200000018000000a0090000f69300008200000000420e40448101880200000024000000bc0900005c9400006001000000440ee008648101880289039204930594069507960897092c000000e409000094950000c204000000440e800970810188028903920493059406950796089709980a990b9a0c000010000000140a0000269a000018000000000e000010000000280a00002a9a00002400000000420e10100000003c0a00003a9a0000040000000000000010000000500a00002a9a0000020000000000000014000000640a0000189a00004201000000420e30428101002c0000007c0a0000429b0000e401000000420e705a810188028903920493059406950796089709980a990b9a0c9b0d001c000000ac0a0000f69c00005600000000420e304a810188028903920493050024000000cc0a00002c9d00007803000000420e50528101880289039204930594069507960897090014000000f40a00007ca000000e00000000420e1042810100240000000c0b000072a000007e01000000420e80015081018802890392049305940695079608000010000000340b0000c8a10000120000000000000010000000480b0000c6a100001200000000000000140000005c0b0000c4a100000e00000000420e104281010014000000740b0000baa100000e00000000420e1042810100140000008c0b0000b0a100000e00000000420e104281010014000000a40b0000a6a100007000000000420e90014281012c000000bc0b0000fea10000bc01000000420e90015a810188028903920493059406950796089709980a990b9a0c9b0d14000000ec0b00008aa30000b400000000420e104281010014000000040c000026a400003800000000420e4042810100100000001c0c000046a400000a0000000000000014000000300c00003ca40000b600000000420e104281010014000000480c0000daa400003a00000000420e404281010020000000600c0000fca400002001000000420ea0014e810188028903920493059406950720000000840c0000f8a500000001000000420ea0014e81018802890392049305940695071c000000a80c0000d4a600009800000000420e4048810188028903920400000014000000c80c00004ca700000e00000000420e104281010014000000e00c000042a700007200000000420e900142810114000000f80c00009ca700007200000000420e900142810110000000100d0000f6a70000160000000000000018000000240d0000f8a70000a200000000420e40468101880289030014000000400d00007ea800007000000000420e90014281011c000000580d0000d6a800005200000000420e304a810188028903920493050018000000780d000008a900007e00000000420e5046810188028903001c000000940d00006aa900006200000000420e2048810188028903920400000010000000b40d0000aca90000360000000000000010000000c80d0000cea90000300000000000000018000000dc0d0000eaa900004e00000000420e10448101880200000020000000f80d00001caa00008600000000420e504c8101880289039204930594060000001c0000001c0e00007eaa00006800000000420e304a8101880289039204930500180000003c0e0000c6aa00007e00000000420e50468101880289030018000000580e000028ab00005200000000420e20468101880289030018000000740e00005eab00005600000000420e10448101880200000020000000900e000098ab00008201000000420e504e81018802890392049305940695070010000000b40e0000f6ac0000280000000000000010000000c80e00000aad00006200000000420e1018000000dc0e000058ad00006800000000420e30448101880200000014000000f80e0000a4ad00003000000000420e104281010024000000100f0000bcad00006601000000420e80015281018802890392049305940695079608970918000000380f0000faae00006400000000420e30448101880200000018000000540f000042af00007800000000420e40468101880289030018000000700f00009eaf00007e00000000420e4046810188028903001c0000008c0f000000b00000a200000000420e5048810188028903920400000018000000ac0f000082b000007a00000000420e20468101880289030020000000c80f0000e0b00000ba00000000420e504c81018802890392049305940600000010000000ec0f000076b1000010000000000000001c0000000010000072b100008c00000000420e404881018802890392040000001000000020100000deb100004a000000000000001c0000003410000014b200007200000000420e50488101880289039204000000100000005410000066b20000c0000000000e0000140000006810000012b300002800000000420e1042810100140000008010000022b300002800000000420e10428101002c0000009810000032b300001401000000420e6058810188028903920493059406950796089709980a990b9a0c00000010000000c810000016b400006c000000000000002c000000dc1000006eb400007e03000000420ed0035a810188028903920493059406950796089709980a990b9a0c9b0d2c0000000c110000bcb700000603000000420ec0015a810188028903920493059406950796089709980a990b9a0c9b0d2c0000003c11000092ba0000e802000000420ec0015a810188028903920493059406950796089709980a990b9a0c9b0d2c0000006c1100004abd0000d002000000420eb0015a810188028903920493059406950796089709980a990b9a0c9b0d2c0000009c110000eabf0000ae02000000420ea0015a810188028903920493059406950796089709980a990b9a0c9b0d14000000cc11000068c200002800000000420e104281010014000000e411000078c200002800000000420e104281010028000000fc11000088c200002801000000420e6056810188028903920493059406950796089709980a990b00200000002812000084c300006800000000420e404e8101880289039204930594069507002c0000004c120000c8c300000403000000440ea00674810188028903920493059406950796089709980a990b9a0c9b0d100000007c1200009cc6000066000000000e00002c00000090120000eec60000c602000000440ef00474810188028903920493059406950796089709980a990b9a0c9b0d2c000000c012000084c900004602000000420eb0025a810188028903920493059406950796089709980a990b9a0c9b0d2c000000f01200009acb00008e02000000440ef00474810188028903920493059406950796089709980a990b9a0c9b0d2c00000020130000f8cd00000202000000420e90025a810188028903920493059406950796089709980a990b9a0c9b0d2c00000050130000cacf00003629000000440ec0046a810188028903920493059406950796089709980a990b9a0c9b0d1800000080130000d0f800008e00000000420e504681018802890300200000009c13000042f90000cc01000000440ec0045881018802890392049305940600001c000000c0130000eafa0000f600000000440ec004548101880289039204930520000000e0130000c0fb00005402000000440ee0045881018802890392049305940600002800000004140000f0fd00000604000000420ee00156810188028903920493059406950796089709980a990b2c00000030140000ca010100e809000000420ec00158810188028903920493059406950796089709980a990b9a0c00002400000060140000820b01005001000000420e9001528101880289039204930594069507960897092c00000088140000aa0c01000c03000000420ed0015a810188028903920493059406950796089709980a990b9a0c9b0d24000000b8140000860f0100c803000000420ec001508101880289039204930594069507960800001c000000e0140000261301006a00000000420ea00348810188028903920400001800000000150000701301008e00000000420e5046810188028903001c0000001c150000e21301007200000000420e50488101880289039204000000100000003c1500003414010028000000000e00001000000050150000481401001c00000000000000200000006415000050140100da00000000440ed0055881018802890392049305940600002000000088150000061501002a02000000420ec0014c810188028903920493059406000018000000ac1500000c1701003200000000420e10448101880200000028000000c8150000221701001803000000420eb00256810188028903920493059406950796089709980a990b2c000000f41500000e1a01008c03000000420ef0025a810188028903920493059406950796089709980a990b9a0c9b0d2c000000241600006a1d01009003000000420e80035a810188028903920493059406950796089709980a990b9a0c9b0d2c00000054160000ca2001004e04000000420e80035a810188028903920493059406950796089709980a990b9a0c9b0d2000000084160000e82401008601000000420e90014c81018802890392049305940600002c000000a81600004a2601005602000000420ef0015a810188028903920493059406950796089709980a990b9a0c9b0d1c000000d8160000702801009a00000000420e6048810188028903920400000018000000f8160000ea2801007801000000420ea001468101880289032c00000014170000462a01005402000000420ef0015a810188028903920493059406950796089709980a990b9a0c9b0d2c000000441700006a2c01007207000000440ea00674810188028903920493059406950796089709980a990b9a0c9b0d1800000074170000ac3301007400000000440eb0044c8101880289033000000090170000043401004a3a000000440ef00f74810188028903920493059406950796089709980a990b9a0c9b0d420e90110000000002452c00014697100000e78060169308d00573000000011106ec22e826e44ae02a890869833589016385a5021796010003368629898db3b4c502998013048503086097900000e780001dfd1413040405e5f80335890001cd03350900e2604264a264026905611733000067006373e2604264a2640269056182800c6591c50861173300006700c3718280797106f422f026ec4ae84ee4aa8508612dc903b9050183b98500630b09060144aa840de426846387090003340422fd19e39d09fe814419a80334052151c883598521850497300000e780e06c8355a4212285e3f3b9fe850991cc8e09a29903b50922fd1491c403350522fd14edfc11c8814911a022857d1981442a84e31309fa39a8a2700274e2644269a269456182806387090003350522fd19e39d09fe8335052199c92e8497300000e780c066833504212285e5f911a02a842285a2700274e2644269a2694561173300006700a36497300000e780206417d5ffff1305c5209305b00297800000e78020240000097186fea2faa6f6caf2ceeed2ead6e6dae25efe62fa66f66af26eee2a8a0061ae8a55c883348a008811a2852686d68697100000e780e0ef0e75630605402e7b03b50a0083b50a014e7cee7d2af8aee003b58a0083b50a0203b68a0283bb8a012afc2ef032f463090b080359ab212d45138d0a026376a90c13851d006362a90213060003b385cd02da953305c5025a95b306b9413386c60297800100e78080ec03b50a0193050003b385bd02da9588e903b50a0088e103b58a0088e523bc750103350d0088f103358d001b04190088f5231d8b20a5a603b50a0183b50a00aae02ef803b58a0083b50a0203b68a0283bb8a012afc2ef032f497000000e78000528355a5212d4663ffc5381b861500231dc520130600038666b385c5024276aa9594e9e27690e10276227794e523bc750190f198f52330aa0023340a00054511a622e405491545914c26e863eead006389ad000149994c63979d01814d954c21a0ee8c11a0e51d97000000e780204b8359ab212a8493c4fcffce94231d952013050003b385ac02da9588111306000397800100e7804098314563f6a42c13851c00b385a9406397953013060003b305c502da953386c402228597800100e780a095231d9b2108198c111306000397800100e7806094da8463130900a28452ec03d9a42113851d006362a90213060003b385cd02a6953305c5022695b306b9413386c60297800100e780e0d503b50a0193050003130a0003b385bd02a69588e903b50a0088e103b58a0088e523bc750103350d0088f103358d00052988f5239d242188080c191306000397800100e780a08c03350b216303051481449549a28a835c8b212a8b08018c081306000397800100e780608a631b9c1e835dab212d4563e6ad1a0549114d63ee3c01668d638b3c01014919456395ac00814c154d19a0e51c194d97000000e780603a8359ab212a849344fdffce94231d9520b3054d03da9588111306000397800100e780c084314563faa418930b1d0033857941631e951813050003b385ab02da95130a00033386a402228597800100e780e081231dab2108198c111306000397800100e780a0808359a42113851900b14563f4b9163386ad416316a616050c8e0bda9b93850b22930404220e06268597700100e780a07d014593153500a6958c6133363501239ca5203295b3b6a90093c61600758e23b8852065f288080c191306000397700100e780607a5a856313090022851001e685d68697000000e780a01b03350b21a28ae2849549e31505ec11a0014c97000000e780c02aaa840355a5218145226623b0c42213890422139635004a961062b3b6a500231cb620b6953337b50013471700f98e23389620e5f2c26513851500626a23309a002334aa00639a850d83d9a4212945636c350d1b851900239da420130500033385a90226958c081306000397700100e78040708509139539004a9500e123389420231c342111a810015a85e685d68697000000e780a010626a03350a0105052338aa00f6705674b6741679f669566ab66a166bf27b527cb27c127df26d19618280ad45268531a817d5ffff130535f19305500315a017d5ffff1305d5ed19a8b14597800000e7808065000017d5ffff130575ec9305800297800000e780e0d9000017d5ffff130525d193050002edb717d5ffff130535eaf1bf17d5ffff130585e493050003c9bf17d5ffff1305c5cee9bf83b605219dc683d78521130816009dc71387f7ff93173700b69783b707222330050014e52338050118ed1cf110f50cf92da00ce510e989450ce1828003d7a62119cf03b7862285471ce114e523380501233c05000cf110f518f910fd828097800000e78020ed00001d7186eca2e8a6e4cae04efc52f856f45af05eec62e866e42a84835aa5213689b2892e8a93841500338bba4063e09a0213060003b305ca02a2953385c40222953306cb0297800100e780009e938b1a00130500033305aa02229513060003ce8597700100e780605793892a00130c042213052a00939c3400637c3501b3059c010e05629513163b0097800100e780c099669c23302c01231d742163f434030e0a229a13058a22b305504109461461239c9620850423b88620b38695002105e397c6fee6604664a6640669e279427aa27a027be26b426ca26c25618280411106e413050022c14597300000e780a0ff01c923380520231d0520a260410182801305002297300000e780e0ff0000411106e413050028c14597300000e780a0fc01c923380520231d0520a260410182801305002897300000e780e0fc0000757106e522e1a6fccaf8cef4d2f0d6ecdae8dee4e2e066fc6af8aa8a0075035ca421330bbc002d45636b65112e8983bb8a0183d4ab2163ebb410338a2441239d4b21231d6421130d00033305a90322953306ac03a28597800100e7802089930c1a00338594419305f9ff6318b50eb385ac03de95b309a50322854e8697700100e780e04103b50a0183b40a00330aaa035e9a3305a503aa940a8513060003a68597700100e780a03f130600032685d28597800100e7808083330534018a851306000397700100e780803d83b50a0203b50a03b9c541c9930404220e093385240113163c002106a68597800100e78000808e0ce69b93850b2226854a8697700100e780e0390145050b8c601306150023b88520239ca520a1043285e317cbfe11a031e1aa600a64e6744679a679067ae66a466ba66b066ce27c427d4961828017d5ffff130575c1930530031da017d5ffff1305c5c39305700221a817d5ffff130535b829a017d5ffff1305b5c49305800297800000e78000a50000357106ed22e926e54ae1cefcd2f8d6f4daf0deece2e8e6e4eae06efc2a89033b8501035cab212e8de2952d456363b5148339890203d5a9216364a515b30ca541231dbb20239d9921930bfdff930d00030335090103340900338abb03ae84b38a49013305b5032a940a8513060003a28597700100e780002b130600032285d685a68a97700100e780c06e3305bc035a958a851306000397700100e780a02893041c0033859a406392ab0e3385b4035a95ce85528697700100e780c026b305bd03ce953386bc034e8597700100e780606a8335090203350903adcd4dcd13840922139534005a951305052213193d00a2854a8697700100e780e022b305240113963c002106228597700100e780806663705c030e0c5a9c13058c220c61239c9520850423b865217d1d2105e3180dfe7d556382ac020145938b1c000c601306150023b83521239ca52021043285e397cbfe11a029e1ea604a64aa640a69e679467aa67a067be66b466ca66c066de27d0d61828017d5ffff1305b5ae930520030da017d5ffff1305f5b011a817d5ffff1305959d29a017d5ffff130515aa9305800297800000e780608a0000557186e5a2e126fd4af94ef552f156ed5ae95ee562e1e6fceaf8eef483bd850103dcad21628701c698750357a7216367d71632ec36f02af483ba850283dcaa21130b1c0033069b012d456360c516806188652ae488712ae883bb05010359a42132e0239dcd20130a0003b3844b03a294081813060003a68597700100e780e00f93891b009385040313c5fbff330d250133064d03268597700100e780e05233054c036e950c181306000397700100e780c00c33054b036e9533864c03d68597700100e780800b93050422139539002e9593943b00a695c10513163d0097700100e780804e63f02903a294138584220c611386190023b88520239c35212105b289e317c9fe0315a4217d358545231da420226563f3a50413153b006e951305052293850a2213963c00210697700100e780c00402656372ac02850c0e0c6e9c13058c22da851061231cb62085052338b621fd1c2105e3980cfe626513341500568597300000e78080b27d143375640182752e95a27523b0b501426690e588e9ae600e64ea744a79aa790a7aea6a4a6baa6b0a6ce67c467da67d6961828017d5ffff130515979305100939a017d5ffff1305459f9305a00297700000e780606e0000717106f522f126ed4ae94ee552e1d6fcdaf8def4e2f0e6eceae8eee4033a850183398502035baa2183dba92113041b0033067401ad4563ebc512833c05000c652ee4833d050103ddac2132e0231dca2013090003b38a2d03e69a080813060003d68597700100e78040f593841d0093850a0313c5fdff330ca50133062c03568597700100e780403833052b0352950c081306000397700100e78020f233052403529533862b03ce8597700100e780e0f093850c22139534002e95939a3d00d695c10513163c0097700100e780e03363f0a403e69a13858a220c611386140023b89521239c95202105b284e317cdfe0395ac217d358545239dac20a26463f29504131534005295130505229385092213963b00210697700100e78020ea02656371ab02850b0e0b529b13058b220c61239c8520050423b84521fd1b2105e3980bfe4e8597300000e78060986685a685aa700a74ea644a69aa690a6ae67a467ba67b067ce66c466da66d4d61828017d5ffff130525879305a00297700000e78040560000457186e7a2e326ff4afb4ef752f356ef5aeb5ee762e3e6feeafaeef6ae8483bb050003ba05013289aa8983daab21130b000333046a035e940a8513060003a28597700100e78040df930504031345faff569533066503228597700100e780a022fd3a13950a03239d5b2183ba8400419195456372b51a2819de85568697f0ffffe780a0776a7505cd85456317b5068001080113068003a28597700100e780c0d96a65aa750355a52183d5a5212e950505b1456376b50408180c01014605a88001a80013068003a28597700100e780c0d60675c6750355a52183d5a5212e950505b145637fb5020818ac000546d28697000000e78000bd89a80e65ae6599a0081a13068003a28597700100e780e0d2081a854597000000e78020a03665d66515a0050a081a13068003a28597700100e780a0d0081a854597000000e7804086766596752af82efcd2e0c27be27a03b60b21066a71c293841a00130b010c914d314c954c054d0354a62163e78d0a2819b285268697f0ffffe78040686a750dcd6318a509a81913068003da8597700100e780a0ca526592750355a52183d5a5212e950505636c8503b3858c40a81997000000e780809691a8a81913068003da8597700100e78060c7526592750355a52183d5a5212e95050563728503081a13068003da8597700100e78020c5081a97000000e78020c92a86ae8409a8b3858c40a81997f0ffffe780a079014629fe29a001e405452300a9008a85130600034e8597700100e78060c123b8790323bc590323b04905be601e64fa745a79ba791a7afa6a5a6bba6b1a6cf67c567db67d796182801d7186eca2e8a6e4cae04efc52f856f45af05eec62e866e46ae0b289ae8a2a89938c0601130a0003854b130bf00f03dcaa21b3044c037d54568595cc130d050341055146e68597700100e78060fc932505003335a000b305b040c98d938404fd05046a85e38b75fd13f5f50f631e65016396090089a06284638f09020e045694833a0422fd1965b701452334590123383901233c89002330a900e6604664a6640669e279427aa27a027be26b426ca26c026d256182802334590123380900233c89000545c9bf130101812334117e2330817e233c917c2338217d2334317d2330417d233c517b2338617b2334717b2330817b233c91792338a1792334b1796d71178601001306e6260ce208e61305014997600000e7802060033501497dc98335014a2d466364b6006f10e002138645ff8d4663e4c6006f1040020346d5008346c5000347e5008347f5002206558e4207e207d98f83461500034705008344250003043500a206d98ec2046204458c03388149c18e91445d8e638c960283465500834745008344650003047500a206dd8ec2046204458cc18e8d47e3f5d716f19ac1476397f60063f4c50432856f00507c938605ff8d4763e4d7006f00b07a83461501834705018344250103043501a206dd8ec2046204458c558c931604029b0706008192e362f478e3e3d578b685918d9146e3e7d576f1159306000263fad502154499446306080097200000e780e04e39a08334014a0334814913d58400220593f5f40f4d8d23388148233ca148cda22a968345c6008346b6008347d6008344e600a205d58dc207e204c58fdd8d834606018347f6008344160103442601a206dd8ec2046204458cc18e821633e4b60083454601834636018347560183446601a205d58dc207e204c58f83468601b3e8b7008347760183449601a2060307a600b3e2f600c2048347a6012303e1340307960083458600e207c58f2207d98d2312b13483455600034746008344660083067600a205d98dc204e206c58ed58d2320b13483053602b3e65700821633e91601230cb1388345c6018346b6010347d6018347e601a205d58d4207e207834606025d8fd98d0347f601a2068347160203462602d98e93548900c20762065d8e558e0216d18d2338b1386306080097200000e780a03b0305613483154134032601342303a12e2312b12e2320c12e1305712f0c0f254697700100e7800088135584032307a12e13550403a306a12e135584022306a12e13550402a305a12e135584012305a12e13550401a304a12e135584002304a12ea303812e13d50403230ba12e13d58402a30aa12e13d50402230aa12e13d58401a309a12e13d504012309a12e13d58400a308a12e2308912ea307212f8544e21493851400054597700000e78020801549114409e993852400054597600000e780e07e29cd23382149233c81481305014997f00000e780e0d1aa8413958403619551618330817e0334017e8334817d0339017d8339817c033a017c833a817b033b017b833b817a033c017a833c8179033d0179833d81781301017f82800545621593051500014597600000e780207845c51305014997600000e780a029833d0149638c0d30833c81490336014a13050149ee8597f00000e78080cb13050002814597800000e780c0ab2a8c2e89930501491306000297600100e780c0729305000205460544628597000100e780c0e31375f50f6300052e130501491306004093040040814597600100e780e0622338913805659b08a5811317840305070c0f130501490146814681470148730000006304052ac94429a32334014a2330014a233c014823380148130500022330a13405659b08e5808c061305014989440146814601478147014873000000630295262a840545630ca4241149e31604ea03340134130500020949e36f85e8032501498315414903066149014d2320a1262312b1262303c1260345814983457149034691498346a14922054d8d4206e206558e518d8345c1490346b1498346d1490347e149a205d18dc2066207d98ed58d8215b3eaa5000345014a8345f1490346114a8346214a22054d8d4206e206558e518d8345414a0346314a8346514a0347614aa205d18dc2066207d98ed58d8215b3eba5000345814a8345714a0346914a8346a14a22054d8d4206e206558e518d8345c14a0346b14a8346d14a0347e14aa205d18dc2066207d98e0346f14ad58d82154d8d2300c132233ca130930d1149130c814a1309713a130b11499309814a130a1139fd5c130501490946ea8597600000e78020ec03450149631f053203856d0083855d0003c64d00230ba138a205d18d231ab13803c51d0083c50d0003c62d0083863d0022054d8d4206e206558e518d0334814983158c0003360c008334014a2328a1382314b1342330c1348c0629464a8597600100e780005113558403230fa13813550403a30ea13813558402230ea13813550402a30da13813558401230da13813550401a30ca13813558400230ca138a30b813813d584032303a13a13d50403a302a13a13d584022302a13a13d50402a301a13a13d584012301a13a13d50401a300a13a13d584002300a13aa30f91388c141d465a8597600100e780a048233c51492330714b2c0e25464e8597600100e78040470345013901cd130600025285da8597700100e78060880125630b0512630e9d41050df1b5033581498335014a97f00000e780609685b9014911a0054991b98144ada4833a01391305104063e7aa068545054a568597700000e7804079aa892e84930501491306004097600100e780404093840ac0138509402338913885659b88a58113178a0305070c0f1306004081468147014873000000833501393335a000b3b5b4004d8d31c9e30b04ce4e8597200000e78000ede5b15685814597700000e780c072aa892e8493050149568697600100e780e039914463f19a0222f54545c54b814597700000e78040702a842e8b17b5ffff9305a55899a003c5190083c5090003c6290083c6390022054d8d4206e206558eb364a60022f563989a12a14463f49a1a4545c54b814597700000e780e06b2a842e8b17b5ffff930545544546228597600100e780a032054d1da21305014997600000e780c0a283340149edc0033a81490339014a1305014d13060004814597600100e780c022130541499309014c1306c002814597600100e780602117b5ffff9305f57341464e8597600100e780002d370501011b0505022328a14823340160080f9305014997400000e7804031080fa6854a8697600100e780800e2338a149080f93050149214697600100e780400d233c0134233801342334013423300134130501490c0f1306800f97600100e780e026130501498c061306000297600100e780600b88068c151306000297600100e780406701257dc963070a00268597200000e780c0d41544154989bc033981490334014aa1b44545c54b814597700000e78080592a842e8b17b5ffff9305e5414546228597600100e7804020014d2328a149232a4149233c91482330514b2334814a2338614b233c714b1305014997600000e780608bc9442a7511c54e8597200000e780c0cd63070900628597200000e780e0cce3870c9e6e8597200000e78000ccc5b203c5590083c5490003c6690083c6790022054d8d4206e206558eb364a60013b5840093f53400b335b0004d8d15cd45454544814597700000e780c04eaa84ae8a17b5ffff930525374546268597600100e78080150d4d91bfe30e0a9c268597200000e78080c5f9b263f09a024545c54b814597700000e780e04a2a842e8b17b5ffff93054533c5bb13d524009305f5ff0d4563f0a5044545c54bae8a814597700000e78020482a842e8b17b5ffff930585304546228597600100e780e00e114d8d44e5b517b5ffff1305252b930510026da02ef16398a50a114611444e85d685a68697500000e780e01b13f63500f199b306b5002338a148233cb1482330d14a2334c14a2338814a080f9305014997500000e78000f2080fd68597500000e780801a033401398334013a23388148233c914809452330a14a1305014997500000e780c02b3dc545454544814597700000e780403daa84ae8a17b5ffff9305a5254546268597600100e78000040d4d69aa17b5ffff1305652ef14597600000e780007500004545c54b814597700000e78060392a842e8b17b5ffff9305c5214546228597600100e78020008d44114d8a7aedbbe38504060545e385a406106014644e85d68597500000e780c00d85c12a86ae8613050149b285368697500000e7802012032d014915456314ad100945e38da402106414684e85d68597500000e780600a85c12a86ae8613050149b285368697500000e780c00e032d014915456319ad0c0d45e388a4001068146c4e85d68597500000e780000785c12a86ae8613050149b285368697500000e780600b032d01491545631ead080335813911c5228597200000e78060a593858aff0d456379b54a93854aff6375b54a03c5990083c5890003c6a90083c6b90022054d8d4206e206558eb366a60003c5d90083c5c90003c6e90003c7f90022054d8d42066207598e3367a60013050149ce85568697500000e78060f7833b014a638a0b04833401495e85814597700000e780a0242a842e8aa6855e8697600100e780e0eb0da8032a414983348149833a014a0334814a033b014b833b814b03358139e30f05c80335013997200000e780209a79b101440335814919c50335014997200000e780c098a944e30004ca0d45636475016f10b0010345140083450400034624008306340022054d8d4206e206558e518d85456314b50a13050149a2855e8697500000e7802019033b01498334014a2685814597700000e780001a2a8dae8bda85268697600100e78040e199e06f10607c034b0d0063870b006a8597200000e780e0900335814919c50335014997200000e780c08f63070a00228597200000e780e08e0545054a6303ab000d4a62151306150013050149814597500000e780a070034501491dc1033581498335014a97e00000e780e02caa84f9b6e3060abc228597200000e780808a7dbe031561498315414903562149834611492312a10ec205d18d033481490335814a0356014b8334014aaed1aae9231cc10c6389062e0315410e8e55231aa10a2ed91305610c8c09294697600100e78040d413550403231ea10a13550402231da10a13550401231ca10a231b810a13d504032312a10c13d504022311a10c13d504012310a10c231f910a130501490c19054697000100e780c0a0033401496305042883048149930591491305110f3d4697600100e780e0cda2f52308910e0802ac1197200000e78060c25265930500026304b5006f102069126583451500034605008346250003473500a205d18dc2066207d98ed58d034655008346450003476500834775002206558e4207e2075d8f598e0216d18d2eee83459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2ef283451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2ef683459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5010345f5012206558e42076205598d518d02154d8d2afa130501492c0a528697f00000e780206b03340149630404148304814993059149130511143d4697600100e78060b922fe2300911463070b120545c944631dab4c13050002814597700000e78020efaa842e8b2c0a1306000297600100e78040b6930500020546054a268597f00000e7804027aa8a63070b00268597100000e780406513f5fa0f930450046316454913050002814597700000e78040eaaa842e8b2c0a1306000297600100e78060b1930500020946268597f00000e7808022aa8a63070b00268597100000e780806013f5fa0f854593046004631fb542228597700000e7806006326511c5126597100000e780205e2e7597700000e780e0042a7511c54e8597100000e780a05c63070900628597100000e780c05b63870c006e8597100000e780e05a81446ff0cfac314521a81145b28509a8114539a0114511a03285b68511a0368597700000e780e0a30000b94461b88344814949b883448149c1a6880a2c1a97100000e780607b080f2c1a97100000e780a06f130501492c1a97100000e7804074033401390336013a833401490337014aa812a285a68697e00000e78020060335814911c5268597100000e78000520335813911c5228597100000e7800051080f2c1a97100000e780205f130501492c1a97100000e780c063033401390336013a833401490337014a2803a285a68697e00000e780a0000335814911c5268597100000e780804c0335813911c5228597100000e780804b28132c1a97100000e7802075080f2c1a97100000e780e04d130501492c1a97100000e7808052033401390336013a833401490337014a8803a285a68697e00000e78060fa0335814911c5268597100000e78040460335813911c5228597100000e780404513050149ce85568697500000e78080f08334014a95c0033b01492685814597700000e78080c9aa8bae8ada85268697600100e780c09011a0814b0335814919c50335014997100000e780804063810b1613050149de85268697500000e780c0c3033b01498334014a2685814597700000e780a0c42a842e8dda85268697600100e780e08b23388138233ca1392330913a88060c0f97700000e78040500335814919c50335014997100000e780603a63870a005e8597100000e7808039033501348335813403360135aaf3aef7b2fba8120c191306000297600100e780c0c801259304600263140518130501490c19054697f00000e780a0550334014961c48304814993059149130511203d4697600100e780e082a2ff23009120130501490c19094697f00000e780805203350149aae845c18304814993059149130591213d4697500100e780a07f46652338a120230c9120a81b97100000e780605f9374f50f080c97100000e780805e1375f50f6393a40e080fac1b97100000e780e071130501490c0c97100000e78000710336013a0335014a6311a604833501490335013997600100e78020bc9334150035a0cd44d9a00145814501bb0545854529b30945894511b38344814955a00d458d45e5b98344814979a081440335814919c50335014997100000e780a0260335813919c50335013997100000e7808025a1cc13050002814597700000e78020ab2a8bae8b2c031306000297500100e78040721305014913060002da8597e00000e78020fb0345014959c18344114963870b005a8597100000e780c020466597700000e78080c701a8466597700000e780c0c693047002228597700000e780e0c51e7597700000e78040c55a7511c53a7597100000e780001d766511c5566597100000e780201c7274228597700000e780c0c2326511c5126597100000e780801a2e7597700000e78040c16ff04fcb03358149aae063870b005a8597100000e7806018280e8c1397100000e78040742330012e2338012e280e97100000e7800066aae46308051e814488062c0e268697100000e780006d130501498c0697100000e780405e0335014ad1456304b5006f1060032330014a0335014983451501034605018346250103073501a205d18dc2066207d98ed58d2320b13a83451500034605008346250003473500a205d18dc2066207d98ed58d034655008346450003476500834775002206558e4207e2075d8f598e0216d18d2338b13883459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f83368149598e0216d18d233cb13889c697100000e78000080c0f51461305014a97500100e780e055080f8c0697100000e780403b8335013a4145e39aa5740335013903448500834b9500834aa500034bb5008345c500aef0034ad500034de5008345f500aeec834505002ee983451500aef483452500aefc83453500aef8834545002ef1834555002ee5834565002eed833581390346750032e189c597100000e78040ff8504a20b33e58b00c20a620bb3655b014d8d220a8675b365ba00420d666662063366a601d18d82154d8da675a2054a66d18d66764206c676e206558ed18d2a6622068a76558eea66c2060a676207d98e558e0216d18d2338b148233ca14888159305014997e0ffffe78040960335013497700000e780209f2665e31d95e08335012f0336812e8336012e03358131233cb1222338c1222334d12297700000e780809c03358120833501207e762338a12e2334b12e2330c12e130501498c1597100000e780e0270335014a93050002e31eb5620335014983459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18d2334b13a83451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2330b13a83459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d233cb13883451500034605008346250003473500a205d18dc2066207d98ed58d034655008346450003476500834775002206558e4207e2075d8f83368149598e0216d18d2338b13889c697100000e78000e10335813a8335013a03368139833601392334a14a2330b14a233cc1482338d14888068c1397100000e780c03f080f866597000100e780c09928140c0f13060149940697000100e780e09f058901e90335012e97700000e780c08221a8ae840335012e13f4f50f97700000e7808081e3160442167593050002e310b54cd66703c5970183c5870103c6a70183c6b70122054d8d4206e206558e518d83c5d70103c6c70183c6e70103c7f701a205d18dc2066207d98ed58d82154d8d2334a14a03c5170183c5070103c6270183c6370122054d8d4206e206558e518d83c5570103c6470183c6670103c77701a205d18dc2066207d98ed58d82154d8d2330a14a03c5970083c5870003c6a70083c6b70022054d8d4206e206558e518d83c5d70003c6c70083c6e70003c7f700a205d18dc2066207d98ed58d82154d8d233ca14803c5170083c5070003c6270083c6370022054d8d4206e206558e518d83c5570003c6470083c667003ee403c77700a205d18dc2066207d98ed58d82154d8d2338a148080f9305014997e00000e780404403340139e30c04000335013a83358139130600053306c5022296233081242334b12432e8233cc124e30f05000665930525002eec33b5a5002af0130504052ae1080f13068003a28597500100e7800012087c2aed6307057c03459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8d233ca1260345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8d2338a12603459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8d2334a1260345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8d2330a1266a652330a12828642c0588e5286088e1080597100000e78080eb8275e390051ce2656366b56a130501498c1497e00000e780c0b90335014a2ae56300056a1306814a086a0c6610622330a12c233cb12a2338c12a2a65233ca12808150ce510e188062c0d97100000e78080eb130501498c0697100000e78000e08335014a4145e390a51a03350149034d8500834a95008344a500034ab5008345c5002efc0344d500034be500834bf50083450500aefc83451500aee483452500aef083453500aeec834545002ef183455500aef8834565002ee98335814903467500b2f489c597100000e78020a4a20a33e5aa01c204620ab3659a004d8d2204e275c18d420be20b33e66b01d18d821533eaa50026652205e6754d8d8675c20566666206d18d4d8dc675a2050a76d18d4a664206a676e206558ed18d8215b3e4a500880697100000e78020ce1374f50f880697100000e780e0d733e644018335013493461400558d3364a6002e8597600000e7800043631b04561c1f03c5170183c5070103c627018386370122054d8d4206e206558e518d232ca12c03c5970083c5870003c6a70083c6b70022054d8d4206e206558e518d83c5d70003c6c70083c6e70003c7f700a205d18dc2066207d98ed58d82154d8d2338a12c03c5170083c5070003c6270083c6370022054d8d4206e206558e518d83c5570003c6470083c6670003c77700a205d18dc2066207d98ed58d8215033481224d8d2334a12c833a812333358000033a0123b305a040b3f555012338a148233c01482330814a2334414b2338a14a233c014a2330814c2334414d2338b14c1305014997700000e780a0c269c9aa84130d0501a8055146ea8597500100e780c01c012571fd03250d01906494608c1d88c903350d0088e103358d0088e536e92330d12e32f12334c12e41cc280e9415a285528697e0ffffe78060180335813149e1033501320336813283350133a30f0132630b06368e052e95033505229305f6ff89c90356a5210e06329503350522fd15edf98355a521fd15233ca136233001382334b13813050149ac1e1306f13397e0ffffe780a0ed8806930501491306000397500100e780c0cf0335014c8336014d8355a52163f9b6322a86a9a602e902f1130501490c0597100000e78080b38335014a4145639ca56c03350149834b850003449500034ba500834ab5008345c5002ef4034ad5008344e500034df50083450500aef4834515002ef883452500aee4834535002efc83454500aefc83455500aef083456500aef88335814903467500b2ec89c597000000e780a077220433657401420be20ab3e56a014d8d220aa275b365ba00c204620d33669d00d18d821533e4a50042752205a6754d8da665c20562766206d18d4d8d8675a2056676d18d46764206e666e206558ed18d8215b3e4a500080597100000e78080a11375f50f85456315b502ca65338595003336b5008a76b3858600b2956385d5000a7633b6c500631f065c014a014da1a84a658a7563e385002685ca652e8a63e39500268a8a75638385002a8a0a752a8d63638500228d4a66333596008a76b38586403385a540058e6306d5008a75b3b5a50021a0ca65b3b5c5009386f5ffb3f5a60033f5c600181f104b146718639307014a90cb94e798e3233cb1482338a14828149305014997d0ffffe78080043365aa01630c0514ba757a768806b405980397f00000e78040aa130501498c06054697e00000e78040a7833b014a63800b48033481491306814a08620c66106a833401492330a12e2334b12e2338c12e10070ce608e2233c7137130501498c06094697e00000e78040a3033b014a63030b44033581499305814a906194659869833501492330c12e2334d12e2338e12e181614e710e3269ab3369a003306a4013696233c613163048600b3368600639e0648b345ba00318d4d8d63100540a81e97100000e780208a1374f50f280e97100000e78040891375f50f9304f0076310a43e8815ac1e97100000e780e08c130501492c0e97100000e780008c0336012f0335014a631da600833501490335012e97500100e780a0e61334150011a001440335814919c50335014997000000e780a0530335812e19c50335012e97000000e7808052630d04365a8597600000e78000f95e8597600000e78060f82a6597600000e780c0f76a6597600000e78020f70a652a84c265e317b58a55a82330a134233401342338b134130501498c061306f13397e0ffffe780c0b825a88335814c0336052111ca835685210357a62185053285e3f7e6fe11a0ae86130500033385a60232958c061306000397500100e78080980345f1339385faff233cb122e30c05c8630b0a3c033504222334a1229305faff2338b12223380520228597000000e78080468db983448139f5a40a640da00a652338a12493041004e1a4834401490a652338a12475ac9304b0035da4426423388124880497d0ffffe78080ca880397e00000e780a04a93751500639505208335812203368123b336b00003370123b307d0407d8e2338d148233c01482330b14a2334e14a2338d14a233c014a2330b14c2334e14c2338c14c233c01301b550501233401321dcd931515002e957d15233ca14c1305014997600000e780a07115c1aa85080f1306000397500100e7808089280e0c0f97d0ffffe780a0d70335814d71f5080f0c0c97000000e780c06d0335013a93050002631fb52a0335013983459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18d233cb13483451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2338b13483459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2334b13483451500034605008346250003473500a205d18dc2066207d98ed58d034655008346450003476500834775002206558e4207e2075d8f83368139598e0216d18d2330b13489c697000000e780e026033581358335013503368134833601342334a13a2330b13a233cc1382338d13888158c1397100000e780e08e8806866597f00000e780a0df280e8c06100f941597f00000e780e0e5058911e9280e97d0ffffe78060b029a89b54850039a0ae84280e97d0ffffe78020af13f5f40f49e5281497d0ffffe78020ae466597600000e78000c61e7597600000e78060c55a7511c53a7597000000e780201d766511c5226597000000e780401c72746fe09fbc8344014905a08344014901a8930400085a8597600000e780a0c15e8597600000e78000c10a652338a1242a6597600000e78000c06a6597600000e78060bf880497d0ffffe780009f281497d0ffffe780a0a546656fe0bff71145de856fe05fbd17a5ffff130585d29305b0026fe0efe01795ffff130565536fe00fe017a5ffff130585d89795ffff938625569305b002901497500000e78080ee00001795ffff1305a5506fe04fdd1795ffff1305e54f6fe08fdc41456fe0bfb717a5ffff1305a5d49795ffff938645509305b00213060149c1b717a5ffff130505d39795ffff9386a55065b717a5ffff1305e5d19795ffff9386854f59bf17a5ffff1305c5d09795ffff9386654e51b717a5ffff1305c5db6fe0afcb97400000e780e057000017330000670083c41733000067004301797106f422f026ec4ae84ee43284ae892a89328597300000e78040c2aa8405c163e38900a2892685ca854e8697400100e78080544a8597300000e78060fd2685a2700274e2644269a26945618280011106ec22e826e42a8497300000e78000beaa8401c926858145228697400100e780c0432685e2604264a2640561828017030000670023f717030000670023f717030000670023f717030000670083fb97000000e78080010000411106e497500000e780a0db0000411106e497500000e780c0da0000397106fc22f82a840a850d4697600000e78060d202650dc14265a26502662af42ef032ec2c08228597600000e780a0fce27042742161828017a5ffff130585bd9795ffff9386253d9305b002300897500000e78080d30000397106fc22f82a840a85114697600000e780e0cc02650dc14265a26502662af42ef032ec2c08228597600000e78020f7e27042742161828017a5ffff130505b89795ffff9386a5379305b002300897500000e78000ce0000397106fc22f82a840a85154697600000e78060c702650dc14265a26502662af42ef032ec2c08228597600000e780a0f1e27042742161828017a5ffff130585b29795ffff938625329305b002300897500000e78080c80000397106fc22f82a840a85194697600000e780e0c102650dc14265a26502662af42ef032ec2c08228597600000e78020ece27042742161828017a5ffff130505ad9795ffff9386a52c9305b002300897500000e78000c30000397106fc22f82a840a851d4697600000e78060bc02650dc14265a26502662af42ef032ec2c08228597600000e780a0e6e27042742161828017a5ffff130585a79795ffff938625279305b002300897500000e78080bd0000397106fc22f82a840a85214697600000e780e0b602650dc14265a26502662af42ef032ec2c08228597600000e78020e1e27042742161828017a5ffff130505a29795ffff9386a5219305b002300897500000e78000b80000397106fc22f82a840a85354697600000e78060b102650dc14265a26502662af42ef032ec2c08228597600000e780a0dbe27042742161828017a5ffff1305859c9795ffff9386251c9305b002300897500000e78080b20000397106fc22f82a840a85394697600000e780e0ab02650dc14265a26502662af42ef032ec2c08228597600000e78020d6e27042742161828017a5ffff130505979795ffff9386a5169305b002300897500000e78000ad0000397106fcaa852800014697600000e78080a6226519cd6265c26522662af82ef432f0081097600000e78000c9e2702161828017a5ffff1305e5919795ffff938685119305b002101097500000e780e0a70000397106fc22f82a840a85054697600000e78040a102650dc14265a26502662af42ef032ec2c08228597600000e78080cbe27042742161828017a5ffff1305658c9795ffff9386050c9305b002300897500000e78060a20000397106fcaa852800094697600000e780e09b226519cd6265c26522662af82ef432f0081097600000e780e0b6e2702161828017a5ffff130545879795ffff9386e5069305b002101097500000e780409d0000797106f422f02a840a85194697600000e780a096026519c94265a265026608e80ce410e0a27002744561828017a5ffff130585829795ffff938625029305b0021306f10197500000e78060980000397106fc22f82a840a85094697600000e780c09102650dc14265a26502662af42ef032ec2c08228597600000e78000bce2704274216182801795ffff1305e57c9795ffff938685fc9305b002300897500000e780e0920000397106fc22f82a840a85014697600000e780408c02650dc14265a26502662af42ef032ec2c08228597600000e78080b6e2704274216182801795ffff130565779795ffff938605f79305b002300897500000e780608d0000797106f422f026ec0c6911466394c500814491a0006110600865050610e031c21306450022e06360a6040d4532e46371b504f1152ee80a8597500000e78060740a8597600000e7806080aa84228597500000e78000532685a2700274e26445618280000000001795ffff1305456729a01795ffff1305a5669305b00297400000e780006a0000797106f422f02a840a8597500000e780807e026519c94265a265026608e80ce410e0a2700274456182801795ffff1305656a9795ffff938605ea9305b0021306f10197500000e78040800000797106f422f02a840a85014697500000e780a079026519c94265a265026608e80ce410e0a2700274456182801795ffff130585659795ffff938625e59305b0021306f10197400000e780607b00001d7186eca2e82a842818054697500000e780c074627539c12665866562762aec2ee832e408102c0097600000e7806089027529c14275a2750276aae4aee032fc2c18228597600000e780409d2265e66046642561175300006700a3401795ffff1305a55d9795ffff938645dd9305b002101021a81795ffff1305255c9795ffff9386c5db9305b002301897400000e780207200001d7186eca2e82a842818094697500000e780806b627539c12665866562762aec2ee832e408102c0097600000e7802080027529c14275a2750276aae4aee032fc2c18228597600000e78000942265e6604664256117530000670063371795ffff130565549795ffff938605d49305b002101021a81795ffff1305e5529795ffff938685d29305b002301897400000e780e0680000057186efa2eba6e7cae3ae842a899385050828001306800f97400100e78060d99385040408021306000497400100e78040d803b4841739cc038504001b05f5fb1375f50f1335050c9335140493c515004d8d39e52800a68597000000e780400613060008018e88022295814597400100e78040c788020c02228697400100e78040d328008c021306000897000000e780c00c39a02800a68597000000e78040022c001306800f4a8597400100e78060d0fe605e64be641e693d618280011106ec22e826e44ae02e892a84130505041306800b814597400100e780c0c01795ffff930545c713060004228597400100e78040cc13053900a14522868346e5ff0347d5ff8347f5ff83440500a206d98ec207e204c58f0347150083442500dd8e834735000217a214458fc217830445005d8f1c62d98ee214c58ebd8e14e2fd1521062105c5fd0345090068f4e2604264a26402690561828069ce797106f422f026ec4ae84ee452e03284ae842a89687193050008b389a54063f6c9082330090e130a09065295a6854e8697400100e78040070335090493050508033689042330b904133505f81345150032952334a9044a85d28597000000e78000083304344113051008ce94636fa402930900080335090493050508033689042330b904133505f81345150032952334a9044a85a68597000000e7804004130404f893840408e3e789fc0335090e4a9513050506a685228697400100e780c0fe0335090e22952330a90ea2700274e2644269a269026a45618280417186f7a2f3a6efcaebcee7d2e356ff5afb5ef762f366ef6aeb6ee72e892a842801130600082401814597400100e78040a80d0941458345e9ff0346d9ff8346f9ff03470900a205d18dc206620703461900d98e03472900d58d0216834639002217598e03074900c216558ed18d6217d98d8ce07d15a104210955fd280213060004a28597400100e78080af2c603064833204053267b2772a65aae89756010083b42612033884053e972a97a58db98d9754010083b4641193d605028215d58d338e9500b346fe004a652ae193d78601a216dd8e2a973303d700b345b30013d70501c215b3e8e500469eb345de0093d6f50386055267d274ea67bee4175501000335250db3ebd50026973e97318d398d9755010083b5650c135605020215518daa95ad8c8a7636f813d68401a214d18c3386e600330996003345a900935605014215b36cd500338abc0033459a009355f5030605f26672772a769754010083b44408b369b500ba96b296328c32f433c59200358d9754010083b424079357050202155d8daa94258fca752eec935787012217d98fae96b382f60033c5a200935605014215b36dd500ee94a58f13d5f703860792761666ea75aefc175701000337470333eba700b296ae963345e800358d17570100033767029355050202154d8d2a97398e8e67bef0935586012216d18dbe96b383b60033c5a300135605014215518d2a97b98dae6a13d6f5038605d18d56934e933345a300135605020215498eb29433c53401ce69935685012215c98e338569004ee8b30ed50033c6ce00935706014216336df600b3009d0033c6d0006e6f9356f6030606b36fd6007a99fae033032b01b347130193d407028217c58f3e97b34467010e75aaf493d88401a21433e61401b3086500b298b3c7f80093d40701c21733e39700330be3003346cb002e75aaf81357f6030606b364e600aa92ae9233c69201135706020216598e329eb345be004e7913d78501a2154d8fb30559004af03388e5003346c800935206014216b36256003386c201318fee751355f7030607336ea700ae93ae86aeecde9333c5b301935d050202153365b501b30c4501b3cd7c01926793d58d01a21db3e5bd00be933e873efcb38db30033c5ad00935305014215336a750033059a01a98d93d7f5038605dd8db69eae9eb3c76e0093d607028217dd8e3696b18d93d78501a215dd8db387ee01b38eb700b3c6de0093d70601c216b3e3f6003383c300b345b30013d6f5038605b3ecc500e298fe98b3c5120113d605028215d18d2e953346f501935686012216d18e56e4338658013696b18d93d70501c215b3e8f500b382a80033c5d2009355f50306054d8d4e982698b3450a0193d605028215cd8eb690b3c5900093d78501a215cd8fb3050701b38ff500b3c6df0093d40601c21633e89600c290b3c6f00093d7f6038606d58fca9df29db3c6ad0193d406028216d58c338f6401b346cf0113d78601a216558fe676ee96338ae600b3449a0093d50401c214c58d2e9f3347ef009354f7030607d98c8a66b69eaa9eb3c5be0013d705028215d98d33871500398d935685012215c98e467b33856e01b30ed500b3c5be0013d50501c215b3eba500338deb00b346dd0013d5f6038606b3e0a600466c62963e96334576009355050202154d8d2a9fb345ff0093d68501a215d58d266e7296b309b60033c5a900935605014215558d2a9fb345bf0093d6f5038605b3edd5002676b29fa69fb3c51f0193d605028215cd8e3693b345930093d48501a215cd8c8675fe95b3839500b3c6d30093d70601c216d58f3e93b346930093d4f6038606b3e8960062673a9a669ab3460a0193d406028216c58eb692b3c4920193d58401a214c58d4279b3044901b38fb400b3c6df0093d40601c21633ea9600b3045a00a58d93d6f5038605d58db29eae9e33c5ae00935605020215c98eb382660033c5b200935585012215c98d33855e01b30cb500b3c6dc0013d50601c216b3eea600f69233c5b2009355f50306053363b50033063b010696b18f13d5070282175d8d3388a400b345180093d68501a215d58d62962e96318d935605014215b360d50006983345b8009355f50306054d8dba93ee93b3457a0093d605028215cd8eb387a601b3c5b70113d78501a215b3e4e500b385c301338a9500b346da0013d70601c216b3e3e6009e97bd8c93d6f4038604c58ee275ae9fc69fb3c47f0113d704028214458f3a9fb3441f0193d58401a214c58d827bde9fae9f33c7ef00935407014217458f3a9fb345bf0093d4f503860533ec95008665ae9caa9c33c7ec00935407020217458fba973d8d935485012215c98ce669338599012695298f935807014217336b1701b30cfb0033c79c009357f7030607b36df700ca8a4a96b305d60033c7be009357070202175d8fb307ef00bd8e93d48601a216c58e66762e96338dc6003346ed00135706014216b36ee600338efe00b346de0013d7f603860633efe6000676329a629a33471a00935407020217458fba92b3c5820193d48501a215cd8c8a68b3854801338a95003347ea00935707014217336cf700e292b3c7920093d4f7038607b3e097004267ba9f9a9fb3c77f0093d407028217c58f3e98b344680093d68401a214c58e2279ca9fb69fb3c7ff0093d50701c217dd8db3870501bd8e93d4f6038606c58e329536953346d501935406020216458e33085600b346d80093d48601a216c58e3a953695298e935406014216336396001a983346d8009356f6030606b362d600569d6e9d3346ac01935606020216d18eb69733c6b701135786012216598e3387a801b30ac700b3c6da0093d40601c216b3e39600b38df30033c6cd009356f6030606558e5e9a7a9ab3c5450193d605028215cd8eb3889601b3c5e80193d78501a215cd8fc675d295338ab700b346da0093d40601c21633ef9600fa98b3c7f80093d4f7038607c58fa675ae9f869fb3c66f0193d406028216d58cb38ec401b3c61e0093d58601a216d58db3863f01b38fb600b3c49f0093d60401c214c58eb69eb3c5be0093d4f5038605c58da66b5e953307c500b98e93d406028216c58eb69833c6c800935486012216458e66753a953295a98e93d40601c21633ec9600b30c1c0133c6cc009356f6030606336ed600e26833871a013e9733466700935606020216558e3303d601b346f30093d78601a216dd8e866a5697330dd7003346cd00135706014216598e3293b346d30013d7f6038606b3e0e600ca894a9a2e9ab3467a0013d706028216d98e3698b345b80013d78501a215d98dc66433079a00b38ee500b3c6de0093d70601c216dd8e3698b345b80093d7f5038605b3e3f5006279ca9f969fb3c5ef0193d705028215cd8fbe9db3c55d0013d78501a2154d8f226bb305fb01338fe500b347ff0093d50701c217dd8dae9d33c7ed009357f70306075d8fc2673e953a95298e9357060202165d8e32983347e8009357870122175d8f2695b307e5003d8e135506014216b362a60016983345e8001356f5030605518d2ae8469d729d33c5a601135605020215498eb29d33c5cd01935685012215c98e06756a95330dd5003346cd00135706014216b36fe600338ebf013346de009356f6030606d18ede9e869eb3c5d50113d605028215d18db388950133c61800135786012216598e33873e01b30dc700b3c5bd0093d40501c215b3ee9500f698b3c5c80013d6f50386054d8e569f1e9fb3458f0193d405028215cd8c2693b345730013d58501a2154d8db3052f01b383a500b3c4930093d50401c214c58db3846500258d1357f5030605498f6665aa97b697bd8d13d5050282154d8daa98b3c5d80093d68501a215d58d8a66be96b380b60033c5a000935705014215336af500b30b1a0133c5bb009355f50306053363b50026794a9d329d33c5a201935505020215c98db388b40033c5c800135685012215498e467c33058d01330fc500b345bf0093d70501c215cd8fbe98b3c5c80013d6f5038605b3e2c500667dea9dba9db3c5fd0113d605028215d18d2e983346e800135786012216518f33866d01da89b30ce600b3c5bc0093d40501c215c58d2e983347e8009354f7030607b36f9700c27dee934265aa9333c7d301935407020217d98cb38ac40133c7aa00135587012217598d027e33077e00b30ea700b3c49e0013d60401c214d18c33865401318d9356f5030605558da666b690aa90b3c6f00093d706028216dd8eb38a060133c5aa009357850122155d8db3878001aa97bd8e13d70601c21633e8e600c29a33c5aa009356f5030605b363d5006a9f1a9f33c5e501935505020215c98d2e9633456600935685012215c98e06657a95330dd500b345bd0013d70501c21533e3e500330fc300b345df0013d6f5038605d18d4665aa9c969c33c69401935606020216558eb29bb3c65b0013d78601a216558fb3862c013309d7003346c900935406014216336b9600da9b33c6eb001357f6030606598ece9efe9e33c74e01935407020217d98ca69833c7f801935687012217d98e3387be01330cd700b3449c0013d70401c214458fb3041701a58e13d5f6038606c98e2275aa97ae973d8f135507020217598db30f7501b3c5bf0013d78501a215d98df297338ab7003345aa00135705014215b362e500969f33c5bf008e689355f5030605b369b500469d329d33450d019355050202154d8db30e950033c6ce00ca7d135786012216598eb384ad01338dc4003345ad00135705014215498fba9e33c6ce00926c9357f6030606b36bf60066993699334669009357060202165d8eb29ab3c6da0093d78601a216dd8ee667ca97338ed7003346ce00135506014216518daa9a33c6da009356f60306063369d6008a652e9c1e9c33468b01935606020216d18e369f33467f004e68935786012216d18f33060c01338bc700b346db0013d60601c216558eb306e601b58fae7493d5f7038607dd8dd294ae94258f9357070202175d8f330f5701b3c5e50193d78501a215cd8fb385b401338cb70033478701935407014217336a9700529f33c7e701ca679354f703060733639700ea97ce973d8d135705020215598db303d500b3c6790013d78601a216558fb3869701b30cd70033459501935705014215b369f500ce93334577006e779357f50306055d8d72975e97398e9357060202165d8eb29fb3c7fb014e7e93d48701a217c58f7297338de7003346a601135706014216b36ae600d69f33c6f7012a779357f60306065d8e5a974a97b3c5e20093d705028215cd8fbe9eb345d901ee6693d48501a215cd8cb305d700b382b400b3c7570093d60701c217dd8eb69e33c7d401aa679354f7030607d98ce297aa97bd8e13d706028216d98eb69f3345f501135785012215598dc697330cf500b3c6860113d70601c21633e9e6004ae3ca9f3345f501ea761357f5030605b36be500e696b2963345da00135705020215598d330ad501334646018a7e135786012216598ef696b30dd6003345b501935605014215558d2a9a334646019356f6030606336bd600429d269d33c6a901935606020216558e329fb3c6e401ea6493d58601a216d58db3069d00b38cd50033469601935406014216458e329fb3c5e501ae6493d7f5038605b3e9f500a6929a92b3c55a0093d705028215cd8fbe93b34573008e7493d68501a215cd8eb3859200b38ab600b3c7570193d50701c217dd8db3877500bd8e13d7f6038606d98e629e369e3345c501135705020215598db302e501b3c6560013d78601a216d98e269e338cc60133458501135705014215b363e5009e9233c556009356f5030605336fd5007af6ee98de9833451601135605020215518d3303f50033c66b00ee76135786012216598ec696b30bd60033457501935605014215336ed5007293334566002e769356f5030605558d66965a96b18d93d605028215d58db386f5013347db00ca67935487012217d98c3e96338bc400b3c5650113d60501c215b3efc500fe96b58c93d5f4038604b3ecb400d69ece9eb345d90113d605028215d18d2e9a33c64901935486012216d18c33860e01b38ac400b3c5550113d60501c215d18d2e9a33c64401ca741357f6030606598ee294aa94a58d13d705028215d98dae96358d2a679357850122155d8d2697330de500b3c5a50113d70501c215b3eee50076e3b388de0033451501126c9356f50306053369d500e29be69b33c57301935605020215c98eb383460133c57c002a77935785012215c98f3385eb00338aa700b3c6460113d70601c216558fba93b3c677002e6893d7f6038606b3ebf600429b329bb3466e0193d706028216d58fbe9233465600ea75935686012216558eb306bb00330bd600b3c7670113d50701c2175d8daa92334656006a6e9357f6030606b369f600f29afa9a33c65f01935706020216d18f3e9333466f00ee66935486012216d18c3386da002696b18f93d60701c217dd8e3693b3c7640093d4f7038607c58fea95be952d8f935407020217d98ca69233c75700935787012217d98fe295b38ab700b3c4540193d50401c214b3efb400fe92b3c5570093d7f503ee74860533eff5007af6d294ca94258d935505020215c98d2e9333456900ce67135785012215498f3385f400330ca700b3c5850193d70501c21533eaf5005293b34567000e7793d7f5038605cd8f5a975e97b98e93d506028216d58dae98b3c61b018a7413d58601a216558d2697b304e500a58d93d60501c21533e9d500ca9833451501aa659356f5030605558db295ce9533c6be00935606020216558eb293b3c6790013d78601a216d98ec2953388b60033460601135706014216598eb293b3c676002e7793d5f6038606d58d56973e97398e935606020216558eb298b3c6170193d78601a216d58fb306c701b389d70033463601135706014216b36ee60076e3f69833c617014e779357f6030606336bf60062972a9733c6ef00935706020216d18fbe93334575008e6f135685012215518d3306f701330cc500b3c7870113d70701c2175d8fba93334575004a6e9357f5030605b36af500f294ae9433459a009357050202155d8daa92b3c555002a7a13d68501a215d18dd294b38c950033459501135605014215336dc500ea92b3c555006e6693d6f5038605b3ebd50032987a98b345090193d605028215cd8eb3846600b3459f004a7393d78501a215cd8fb30568003389b700b3c6260193d50601c216d58dae94a58f93d6f7038607dd8e4e963696318f9357070202175d8f33085700b3c60601ea6713d58601a216558d3e96b30dc5003347b701135607014217b369c7004e98334505011356f5032e670605336fc5007af662975a973345ed00135605020215518db302950033465b009357860122165d8e5297330be60033456501135705014215336ae500d292334556001356f5030605518de69fd69fb3c5f50113d605028215d18d3387150133c6ea00ea74935786012216d18f33869f00b38fc700b3c5f50193d40501c215b3e895004697b98f93d5f7038607dd8d4a9e5e9eb3c7ce0193d407028217c58fbe93b3c47b0013d68401a214458e7293b30e6600b3c7d70193d40701c217c58fbe933346760092649356f6030606558eee94aa94a58f93d607028217dd8e3383e600334565000e779357850122155d8d2697b30be500b3c6760193d70601c21633eef60072e3729333456500ce669357f50306053369f500da96ae9633c5d900935705020215c98fbe9333c57500ee75935485012215c98c3385b600338ba400b3c7670193d50701c217dd8dae93b3c674008a7a93d7f6038606b3e9f600d69fb29fb346fa0193d706028216dd8e369833460601ae77935486012216458efe97330cf600b3c6860193d40601c216c58e369833460601ce741355f6030606336aa600a69efa9e33c5d801135605020215518daa9233465f002a67935486012216458eba9e330fd6013345e5019357050142155d8daa92334656009357f60306065d8e5e973297b98d93d705028215dd8d2e9833460601ca67935486012216d18c3306f700b38cc400b3c5950113d70501c215b3efe5007e98b3c5040113d7f503ea678605b3eee50076f6da97ca97bd8e93d506028216cd8eb3885600b345190113d78501a2154d8fb3855701330bb700b3c6660193d70601c216b3eaf600d69833471701aa779354f7030607458fe297ce973d8d935405020215458d2a93b3c46900ca7693d58401a214c58dbe96b38bd500334575019356050142153369d5004a9333c56500ea759356f5030605c98efa95d2953345be00935405020215c98ca69333457a008e67135685012215498e3385f500330ca600b3c4840193d50401c214c58db38775003d8eae629354f6030606458e969cba9cb3c5950193d405028215c58db3836500334777004e63935487012217458fb3846c00330d9700b3c5a50113d50501c21533efa500fa9333457700ee6c9355f5030605b369b500669b369b33c56f019355050202154d8daa97bd8e8e7513d78601a216d98eda95338bb60033456501135705014215498f330ef70033c5c601ae769357f5030605336af500de96b29633c5da009357050202155d8d2a9833460601ce7f935786012216d18f3386f601b38bc70033457501935605014215558d2a98b3c50701ee7793d6f5038605b3ead5003e9c769cb345890193d605028215d58dae98b3c41e01926613d68401a214458eb304dc0033099600b3c5250193d40501c215c58dae98334616019354f6030606458eea97b2973d8f935407020217458f3a9833460601935486012216458ee697330cf60033478701935407014217b36e97007698334606011357f6030606aa74598e7ae332f6da94ce94258d135605020215518d3306150133c7c900935787012217d98f33875400b389e70033453501935405014215b36895004696b2ea3d8e1355f6030606b367a6005e93529333c565009355050202154d8daa93b3457a0013d68501a215d18d3306d3003383c50033456500935605014215b362d500969333c575009355f5030605b366b500ca9fd69f3345ff01935505020215c98d2e9e33c5ca01ea74135685012215498e33859f00330fa600b3c5e50193d40501c215cd8c269eb345c6014a6613d5f5038605c98d62963e96b18c13d504028214458daa93b3c77700ae7413d78701a2175d8f26963a9632e6318d135605014215518d2ae31e95aaee398d1356f5032a670605518d2afa4e97369733c5ee00135605020215518d2a9e33c6c601ea669357860122165d8eba96b29636ea358d935605014215558daaf67295aaf2318d1356f5038e760605518d2afe9a96ae9633c5d800135605020215518d2a98b3c505010e6613d78501a215d98d36962e9632ee318d135605014215518daafa4295aae62d8d9355f50306054d8daae23275ca75aa95fa9533c6b200d666135706020216598eb296358d0a779357850122155d8dba95aa952ef2b18d13d60501c215d18daefeb695aeea2d8d9355f5030605c98da8022ef6a1451060833605fc1861358e398e10e0fd1521052104f5f5be701e74fe645e69be691e6afa7a5a7bba7b1a7cfa6c5a6dba6d7d6182801d7186eca2e8a6e4cae02e89aa840a8513060004814597200100e780a0fae8749305000263e9a50aa86855e5e870ac603386a500b46403c7040fb335b600b0e0b695ace419c3fd55acecfd5513061008ace86378c50813060008138404066309c500098e2295814597200100e78080f52685a28597e0ffffe780e04921459305310026861462a38ed5fe13d78600238fe5fe13d70601a38fe5fe13d786012380e50013d70602a380e50013d786022381e50013d70603a381e500e1922382d5007d152106a1055dfdf0748a854a8597200100e78000fce6604664a6640669256182809305000897300000e78020f70000657106e722e3a6feae842a84938505080a851306800f97200100e78080f8a81913060004a68597200100e78080f793850404281a1306000497200100e78060f683b6841789ca0a85ac19301a97200100e78040d439a00a85ac1997200100e78040c98a851306800f228597200100e78040f3ba601a64f67459618280197186fca2f8a6f4caf0ceecd2e8d6e4dae05efc62f866f46af06eec906103bc8500329c636fcc34aa8988699376f50093b616003337a000f98e6380063a814a89466368d5008d462a87850a0581e3ede6fe83cb85013285d68597000000e780a03b6365ac322a8d1305000463f5aa323305ac4133555501814c89456368b5008d452a86850c0581e3edc5fe938d2c0063ea9d316145b3b5ad02639a0530b384ad02ea9463eaa43113893c006a847d19268a630d0902630c0d24233044015285639b0b00130600105285814597200100e78080d80860610408e1c10408e5e3f844fd1775ffff130525f0a5ac4ee0638b0d2e014b13098d0093891c005a85ee8597000000e780a03563030d201d05935435002330490163990b0052858145268697200100e78040d3d29463e24425638669016109050b268ad1b7094963e72d0593098d02330a904105442285ee8597000000e780c0301d05135b350023b0990063990b00268581455a8697200100e780a0ce33856401636195200504b3058a00e109aa84e39325fd11a02685d68597000000e7806028636fac2463860d262a8b938bfdff2a84638b0b161385edff9305f00363eda520854c5a846ae86ee463080d14aa843395ac00331d55013309a401636589186145b38da402c265ae9d3385ab022e9593098500130a0501636f2c0d03b50d000c612300b40013d68503a303c40013d605032303c40013d68502a302c40013d605022302c40013d68501a301c40013d605012301c400a181a300b40093558503a307b400935505032307b40093558502a306b400935505022306b40093558501a305b400935505012305b40093558500a304b4002304a4000c6180e500e15a85d6852686a28697000000e780c022058915ed5a85d6855e86a28697000000e780802183b5090013563500b295838605001d893395ac00c98e2380d50083350a00b29503860500518d2380a5004a846a99e37489f249a82685a26597000000e780c0185a85d6852686a28697000000e780801c83b58d0013563500b295038605001d893395ac00518d2380a50081cc1385f4ffa68b426de31c0dea97200000e780804f0000426da26d63638c0a33058c40826523b0650123b4850188e923bca50123b0b50323b45503e6704674a6740679e669466aa66a066be27b427ca27c027de26d096182801775ffff1305a5c8f14597200000e780402e00001775ffff130565c7f5b71775ffff1305c5c6cdb71775ffff130525c6e1bf1775ffff130585bfada81775ffff1305e5c193054002c9b71775ffff130505c45dbf1775ffff130565baa1a81775ffff1305c5c24db71775ffff130525bc91a01775ffff130585b59305300271b71775ffff1305a5c429a85285d68597000000e780c002637bac001775ffff130585c797000000e780400500001775ffff1305e5b79305100289bf01cd1306000463f0c5027d153355b50005053315b50082801775ffff130585b59305100239a01775ffff1305a5b79305400297200000e7802020000097200000e780403c000063efa5006382a5021345f5ffaa951305000463f2a50205453315b50082801775ffff1305c5b029a01775ffff130525b09305100239a01775ffff130545a99305300297200000e780c01a000063e0a6041307f003636cc7001307000463fde500898e33d5c6003355b50082801775ffff1305e5ae29a01775ffff130545ae9305400297200000e780c01600001775ffff130565b9b545f5b790659461137806fc3698636bd80c98699355660063e3e500ba8594e2094694e6b68763ebc508fd1593d8860393d2060313d3860293d3060213de860193de060113df8600b68736863e879387070463efe7062380c70013578603a383e700135706032383e70013578602a382e700135706022382e70013578601a381e700135706012381e7002182a380c7002384d700a387170123875700a386670023867700a385c7012385d701a384e70190621ce6fd159ce23e86c9f99385070463e7f50214e1233405010ce914ed82801775ffff130565a2f14597200000e780000800001775ffff130525a1f5b71775ffff130585a0cdb7717106f522f126ed4ae94ee552e1d6fcdaf8def4e2f0e6eceae82a841305000497350100138ae5ff6371850417350100930425ff8860631e05348864fd558ce063130512c870cc6cd068d464aae4aee032fc36f80a850c1897000000e780209c054588e413850401c5a803350a04631b053203358a04fd552330ba041ded03350a0883358a0703360a07aae02efc32f80a850c1897000000e78080e705452334aa040265a2654266e2662338aa04233cba042330ca062334da0603398a0663000902033509000c6110650ce20c6510610ce6130b0a04630825032a8991a403390a0603358a056373a902130509046368252983350a042330aa0685052330ba046315092209a823340a0619ac03350a0405052330aa0403350a00631e052803358a00fd552330ba001ded03350a0a83358a0903360a0983368a08aae4aee032fc36f80a850c1897000000e780408d05452334aa0013050a018a851306000397100100e780e07d83398a031305f003636335210545814c3315350163788500850c63840c1c0605e36c85fe83350a0363e3bc00e68503358a020146e146b386dc02aa96138406fdb385bc406389c516630d051c147803b9060061047d16e307d9fe033509008335890088e1033589008335090088e5047017350100130b85e403350b0183358b03934af6ffe69a5686ca8697000000e78000cd93553500a695038605001d89854b3395ab00518d2380a50063f85c11130c000417350100130b65e0138afaff63778a1333954b01b3143501ca9463e72413033d840203350b0183358b035686ca8697000000e780a0c793553500ea95038605001d893395ab00518d2380a500833a840003350b0183358b035286ca8697000000e780c0c493553500d695038605001d893395ab00518d2380a50008600c612380b40013d68503a383c40013d605032383c40013d68502a382c40013d605022382c40013d68501a381c40013d605012381c400a181a380b40093558503a387b400935505032387b40093558502a386b400935505022386b40093558501a385b400935505012385b40093558500a384b4002384a4000c6184e504e12114d28ae3e54cf119a00149528b03350b0005052330ab004a85aa700a74ea644a69aa690a6ae67a467ba67b067ce66c466d4d6182801765ffff1305656b21a81765ffff1305c55e9305300231a01765ffff1305e569f14597200000e78080cf00001765ffff1305a55cf9bf1765ffff13050568cdb797200000e78080e900001775ffff1305d5a19765ffff9386455815a01775ffff1305b5a09765ffff9386255709a81775ffff1305959f9765ffff93860556c1450a8697200000e78080e40000317106fd22f926f54af14eed52e956e55ae1defce2f8e6f4eaf0eeec97350100938ce5c283b50c04639d05382a8903b58c04fd5523b0bc041de917350100130405c148602c7c3078aae4aee032fc28002c1897000000e78060ae054528e42265c2656266827628e82cec30f034f403b50c0583b58c053335a9001345f5ffb335b9006d8d51c517350100130545bc2c75638e052090612300c90093568603a303d900935606032303d90093568602a302d900935606022302d90093568601a301d900935606012301d9002182a300c90013d68503a307c90013d605032307c90013d68502a306c90013d605022306c90013d68501a305c90013d605012305c90013d68500a304c9002304b900906165a203b50c0483b50c00050523b0ac04639b052a03b58c00fd5523b0bc0015ed173501001304c5b148704c6c50685464aae8aee4b2e036fc28002c1897f0ffffe780c04f054508e4130504012c001306000397100100e780804083ba0c03638f0a2283b98c02138afaff13848902854463809a04638b0922033b040003b50c0183b58c032686ca8697000000e780609593553500da9583c505001d8933d5a50005898504610469d5f91463e6440139a263030a108144930a0004268b63e49a00130b000483bb8c0303bc0c0161453385a4024e9513048502054d03b50c0183b58c032686ca8697000000e780808f638e091a833504fe13563500b2950386050093767500b316dd0093c6f6ff758e2380c500937515003306b040833604fe13661600329513563500369603460600937675003356d600058a51e2630b9b1263fe5b1333159500331575016295636e85131061146590e21065146190e691c12a89833d040003b50c0183b58c0385042686ca8697000000e780c08693553500ee95038605001d893315ad001345f5ff718d2380a5006104e3129af4d28405a023302901930585064a862334260123b02501930c050451a8638a090e814461453385a4024e9508610c612300b90013d68503a303c90013d605032303c90013d68502a302c90013d605022302c90013d68501a301c90013d605012301c900a181a300b90093558503a307b900935505032307b90093558502a306b900935505022306b90093558501a305b900935505012305b90093558500a304b9002304a9000c6123b425012330250103b50c00050523b0ac00ea704a74aa740a79ea694a6aaa6a0a6be67b467ca67c067de66d296182801765ffff1305c51e29a01765ffff1305251e9305300231a01765ffff13054529f14597200000e780e08e00001765ffff1305052293051002edb797200000e78040a900001765ffff130595619765ffff9386051809a81765ffff130575609765ffff9386e516c145300097200000e78060a500005d7186e4a2e026fc4af84ef452f056ec83ba050263800a0a2e8a2a898065b35954034e8597000000e780200b83340a002ae02ee402e863e335078145636e54031396350032950d466370560983c6140003c70400a206d98e03c7240083c7340033045441d6944207e2075d8fd98e14e185052105e37a54fd2ee8226502662338b9002334a9002330c900a6600664e2744279a279027ae26a616182800a8581454e8697000000e7806008c2650265e37954f9d9b71765ffff13054523e54597100000e780e07d00001145d68597200000e78040070000011106ec22e826e42a841dc51355c40305ed93351500931434008e0599c4268597d0ffffe780a0b8aa8581e9268597d0ffffe780c0b90000a1452e85a285e2604264a2640561828097d0ffffe780c0b80000411106e497000000e78000037d567e1605066315c500a2604101828011e597d0ffffe78040b600002e8597d0ffffe780e0b400005d7186e4a2e026fcae86b29563f4d5000145a1a82a8408659314150063e39500ae84914563e39500914493d5c40393b51500139634008e0501c914600e0536f0a14636f42af811a002f42800141097200000e7800028a265426599c1e26531a008e004e47d557e150505a6600664e27461618280411106e4054697000000e78060f87d567e1605066315c500a2604101828011e597d0ffffe780a0ab00002e8597d0ffffe78040aa0000797106f422f026ec4ae84ee452e06365d7046366e604aa89b304d7403389d5002685814597200000e780802c2a842e8aca85268697100100e780c0f323b0890023b4490123b89900a2700274e2644269a269026a456182803685ba8519a03a85b28597200000e78080ed000063e8c60063e9d500b385c640329582803285b68511a0368597200000e78060eb0000011106ec22e826e42a8410690865ae846319a6002285b28597000000e78040f210680860931536002e9504e1050610e8e2604264a26405618280397106fc22f826f44af04eec52e856e4114a32892a84637d46032d45ad4a814597200000e7804020aa84ae891765ffff930505042d46268597100100e78000e7054508c0233444012338240104ecb1a803c5150003c6050083c6250083c535002205518dc206e205d58db3e4a500b9c09104638424052d45ad4a814597200000e780801a2a8aae891765ffff930545fe2d46528597100100e78040e12320040004e423382401233c4401233034032334540331a0114a631d4901154508c0e2704274a2740279e269426aa26a216182802d45ad4a814597200000e780e014aa84ae891765ffff9305a5f82d46268597100100e780a0db23200400a9b71061833805011c65210605483e8763ee17019307f7ff10e11ce5637d1801833686ff0c622106e3f3d5fe333517011345150082800545854597200000e780e0d30000797106f422f026ec4ae84ee452e02e89aa8413050002130a0002814597200000e780a00c2a84ae8913060002ca8597100100e780c0d380e023b4340123b84401a2700274e2644269a269026a45618280397106fc22f826f44af0b2841106636996042e892a843285814597200000e780c0072ae02ee402e826ce10100a856c0897200000e780e0ec330699000a85ca8597200000e780e0eb4265a265026608e80ce410e0e2704274a2740279216182801765ffff1305c5e4f14597100000e780603d0000797106f422f026ec4ae84ee452e08d4663f3c604aa899304c6ff138945002685814597200000e78000002a842e8aca85268697100100e78040c723b0890023b4490123b89900a2700274e2644269a269026a456182801145b28597200000e78060c10000011106ec22e826e44ae02a841305000285451309000297c0ffffe780607329c9aa8413060002814597100100e780c0b404e0233424012338240111458545914497c0ffffe780c0701dc5a301050023010500a30005002300050008ec04f004f423080402e2604264a2640269056182801305000211a0114597c0ffffe780406f0000757106e522e1a6fccaf8cef4d2f0d6ecdae8dee4e2e003bb050193040b0163e86415938b140063890b142e8a83ba8502b3895b0163e779152a894e85814597200000e780e0ef2ae42ee802ec0d4597000000e78020ad2af02ef402f899c1814501a8081097000000e78060bbc27502758e052e95c1450ce1c27585052ef822756398a500081097000000e78040b9c275027c13953500629504e19384150026f82275639aa4000810a68597000000e78000b7c274027c1394340033058c00233075014ede900028006c1897200000e780a0cda2797d556384a402930b0104210462850c61930485002ede28006c185e8697200000e78040cb611426857df063870900628597c0ffffe780e05c83350a0013040a0333866501280097200000e780a0c813061a032800a28597200000e780a0c783358a0133865501280097200000e78080c66265c26522662338a9002334b9002330c900aa600a64e6744679a679067ae66a466ba66b066c496182801765ffff130545be11a81765ffff1305a5bd29a01765ffff130505bdf14597100000e780a01500000d476371c7069306c6ff637ad704930686ff0d476375d70403c8550003c7450083c7650083c6750022083367e800c207e206dd8ed98e03c8950083c8850083c2a50083c7b500220833671801c202e207b3e757005d8f17030000670043a61145b68519a01145b28597200000e780c0980000411106e410610e069766ffff93862681369610620286907588711c6e9765ffff938595c33d4635a8907588711c6e9765ffff9385c5c12d462da021052ae01765ffff9307c5bd1765ffff130745be3d463da0907588711c6e9765ffff9385a5ba2146a2604101828721052ae01765ffff9307b5b61765ffff1307e5b61d468a862e85be8597200000e7806086a2604101828082808365050005466345b60099c9054609a809466389c5000d466394c500210521a0610511a041050c6591c5086117c3ffff6700a3408280130101ba233c1144233881442334914423302145233c3143233841432334514323306143233c71412a8b08081306004013040040814597000100e780a07e2338814005659b0895819305014105470808014681468147014873000000aa84094505446384a412638084081144639f0410033a0141130500406379450785450544528597200000e78080beaa892e890c081306004097100100e780a08593020ac0138509402338514085659b88958193050141130600400547094381468147014873000000630c650aaa846308850a1144d5e483340141094463e2920a13054afd1334150035a001444da05285814597200000e780c0b7aa892e890c08528697000100e780007f1305c00201446306aa023d45bd4b814597200000e78040b5aa84ae8a1765ffff9305b59c3d46268597000100e780007c01c823303b0123342b0123384b0189a802c81305c0022aec52f026f456f85efc0d452334ab0023300b00080897000000e78080e6630609024e8597c0ffffe780002939a80144630709004e8597c0ffffe780e02723348b0023389b0023300b008330814503340145833481440339014483398143033a0143833a8142033b0142833b8141130101468280397106fc22f83287ae862a8402f002ec02e802e4130500022af405659b0815822c108d472800894201460148730000006309550285456308b502914515e522751306000289456361a602130514002c001306000297000100e780a06d2300040009a8854511a081450ce408e805452300a400e270427421618280397106fc22f83287ae862a8402f002ec02e802e4130500022af405659b0815822c109547280089420146014873000000630b55028545630cb502914515e922751306000289456365a602130524002c001306000297000100e780006601458545a300b40009a80145a300040029a081450ce408e805452300a400e270427421618280130101ba233c1144233881442334914423302145233c3143233841432334514323306143233c7141b289ae8b2a8408081306004093040040814597000100e780a0522338914005659b08c58293050141080889440146de864e8781470148730000006301950885456300b508914535ed03390141130500406372250b8545054b4a8597200000e780c0922a8aae8a0c081306004097000100e780e059930209c013050a402338514085659b88c58293050141130600408944de864e87814701487300000063019508630e6507114b25ed03350141094b63e8a2062330440123345401b1a8854511a081450ce408e8233004008330814503340145833481440339014483398143033a0143833a8142033b0142833b81411301014682804a85814597200000e780e088aa84ae890c084a8697000100e780205004e0233434012338240145bf014b2334640108e823300400e3810afa528597c0ffffe780e0fe51bf130101b8233c1146233881462334914623302147233c3145233841452334514523306145233c714323388143233491432330a1432a8d28001306004013040040814597000100e780203c2334814005659b08458093058140280009440146814601478147014873000000aa84630f85060545638ea4061144639b0412833b81401305004063777507854505445e8597100000e780007caa892e892c001306004097000100e780204393820bc0138509402334514085659b884580930581401306004009438146014781470148730000006308650caa846304850c1144f1e083348140094463ee920aa1a00544c9a001447da85e85814597100000e7808075aa892e892c005e8697000100e780c03c114a63f04b033145b14c814597100000e7804073aa8a2e8b1755ffff9305f55925aa03c5190083c5090003c6290083c6390022054d8d4206e206558e336aa60063934b03214a63fe4b093145b14c814597100000e780006faa8a2e8b1755ffff9305b555d5a83145b14c814597100000e780406daa8a2e8b1755ffff9305f5533146568597000100e78000348144e1a80144630709004e8597c0ffffe780e0e323348d0023389d0023300d008330814703340147833481460339014683398145033a0145833a8144033b0144833b8143033c0143833c8142033d014213010148828003c5590083c5490003c6690083c6790022054d8d4206e206558e336aa60013358a0093753a00b335b0004d8d15c53145b14a814597100000e780a0622a8aae8b1755ffff930555493146528597000100e78060298d443da063ff4b053145b14c814597100000e780c05faa8a2e8b1755ffff930575463146568597000100e7808026854426c462c652e85eec56f05af466f80d452334ad0023300d00280097000000e7800092e30209f24e8597c0ffffe78080d419bf13542a007d140d456379a4023145b14c814597100000e7806059aa8a2e8b1755ffff930515403146568597000100e78020209144a28b0d4a59bf6316a408114611444e85de85d28697f0ffffe780002e13f63500f199b306b5002ae42ee836ec32f022f4130581402c0097f0ffffe780c00413058140de8597f0ffffe780202d833a81400334814156e422e809452aec280097f0ffffe780e03e29cd3145b14a814597100000e78060502a8aae8b1755ffff930515373146528597000100e78020178d4411aa3145b14c814597100000e780c04daa8a2e8b1755ffff930575343146568597000100e780801491440d4aa28bf1bd6304041005456304a41003b60a0083b68a004e85de8597f0ffffe780e021130a0002639b450709456306a40e03b68a0083b60a014e85de8597f0ffffe780c01f054a639b45070d456309a40c03b60a0183b68a014e85de8597f0ffffe780c01d2a86ae862800b285368697f0ffffe7806022a24415456392a4080335014111c5568597c0ffffe78080bc23303d0123342d0123387d0169b32e8c3145b14c814597100000e7804041aa8a2e8b1755ffff93054524314605a02e8c2945a94c814597100000e780403faa8a2e8b1755ffff9305a5212946568597000100e78000068144e28b03350141e30905de0335814097c0ffffe780a0b5cdb3324c426ae26b827a227bc27cf9bf0145814509a80545854531a00945894519a00d458d4597100000e78040fe00009308d0057d558145014681460147814701487300000001a041112e87aa8602e405659b0875812c000545014681470148730000001335150041018280086101a08280797106f42e8813564500130f7002130710279756ffff938ee62e6363e608130f700213076102171601008338a66239661b03068f05669b03b6479302c0f937e6f5051b0ef60faa86333515032d813b066502b307d600139607034992330676029355160141821376e67fbb855502be95769683471600c615c19103460600a30ff7fef69583c7150083c50500711f230fc7fea300f7002300b7007117e365defa130630066370a60493150503c99105661b06b647b385c502c5811306c0f93b86c502329546154191791f7695034615000345050093061100fa96a380c6002380a6002e85a945637cb5009305ffff130611002e961b0505032300a60005a006059305efff7695034615000345050093061100ae96a380c6002380a60093061100ae96130770020d8f1755ffff9305855d4285014697000000e780e000a27045618280597186f4a2f0a6eccae8cee4d2e056fc5af85ef462f066ec6ae86ee4aa8403654503ba893689328aae8b937c1500b70a110063840c00930ab00293754500ce9c89e5814b8c6085e5a1a08145630e0a005286de86038706008506132707fc134717007d16ba957df6ae9c8c6095c103bd840063ffac01218925ed83c58403054633059d41634cb60af9e1aa8c2e85c9a0807084742285a6855686de86528797000000e7806014054b0dc15a85a6700674e6644669a669066ae27a427ba27b027ce26c426da26d656182809c6c2285ca854e86a6700674e6644669a669066ae27a427ba27b027ce26c426da26d6561828780581305000383c584032ee003bc040283bd840288d8054b238c64036285ee855686de86528797000000e780e00c51f5228a33049d4105047d1451c803b60d02930500036285029665d985bf09466398c50093051500058193dc150011a0814c03bc040203bd84028458130415007d1409c803360d026285a68502966dd9054b2dbf37051100054be389a4f26285ea855686de86528797000000e780e00511fd83368d016285ca854e86829619f5b30990417d5a7d59338529016309450303360d026285a6850296050975d50da083b68d016285ca854e868296e31005ee014b23a844030265238ca402c1bd6689333b9901e1b5797106f422f026ec4ae84ee49b070600370811003a89b6842e84aa896389070114704e85b2858296aa85054591ed81cc1c6c4e85a6854a86a2700274e2644269a269456182870145a2700274e2644269a269456182805d7186e4a2e026fc4af84ef452f056ec5ae85ee483320500146933e7d2003289ae896304072a638706101c6d8146338e29018507370311009308f00d1308000f4e8601a893051600918eae962e866303640efd17adc7630fc60d8305060013f4f50fe3d105fe834516009374f40113f7f50363fa8802834526001a0793f5f503b363b7006367040383453600f614ad909a0393f5f50333e4b300458c630c64089305460055b79305260013946400598c61bf93053600b20433e4930071b7630bc6078305060063d3050493f5f50f1307000e63ede5021307000f63e9e50203471600834726001377f70393f7f70303463600f615ad9132079a075d8f1376f603598ed18d370611006386c50285c263fd2601b385d90083850500130600fc63d7c500814591e539a0e39d26ffce8599c13689ae89638b021803388500930500026372b902814e63060916ca85ce86038606008506132606fc13461600fd15b29efdf581aa13877900619b3386e940b308c90093f678008145630d3701ce87038407008507132404fc934414000506a6957df6014691ce93f788ffba9783840700850793a404fc93c41400fd162696fdf693d638009717010083b787129714010083b28412b714001092048504939804018508b30eb6001da013173e001a97b386c34113763e00b3f45500a181b3f55500a695b3851503c191ae9e2deaddcab6833a839305000c368e63e4b600130e000c9375ce0f139435001a94dddd81451a8745df146393c4f6ff9d8099821067c58efd8eb6959346f6ff9d82046b1982558e7d8e93c6f4ff9d829980c58e046ffd8e3696b29513c6f4ff1d829980458e7d8e13070702b295e31d87fabdb7630803029305000c63e4b3009303000c814593f633008e06106021041347f6ff1d831982598e7d8ee116b295f5f611a0814533f65500a181b3f55500b295b3851503c191ae9e63fc0e01834685030546b305d8416345d60285ce814a25a80c7508719c6dce854a86a6600664e2744279a279027ae26a426ba26b6161828709466398c600138615008581935a160019a0ae8a8145033b0502833b85020459138415007d1409c803b60b025a85a68502966dd9054a81a037051100054a638ca40283b68b015a85ce854a86829605e533095041fd597d5433058900630a350103b60b025a85a6850296050475d511a05684333a54015285a6600664e2744279a279027ae26a426ba26b61618280411106e497000000e780801c0000197186fca2f8a6f4caf0ceecd2e8d6e4dae0b2891306000232f80d46230cc10203b4090202e002e82af02ef461c003b589026307051083b409009305f5ff8e058d8113891500a10493058003330ab5026104854a17050000130b458a906001caa276027583b584ff946e829665ed08482ad803058401230ca1024c4803b509012eda033684ff0c6001ce631756019205aa95906563046601014621a08c618c61054632e02ee4033684fe833504ff01ce631756019205aa95906563046601014621a08c618c61054632e82eec0c6492052e95106508618a85029649e5c104130a8afc13048403e31b0af6b1a003ba890163080a0483b4090103b409001305faff12051181130915002104a104120a106001caa2760275833584ff946e829639e1906003b584ff8a8502960ded4104411ac104e31e0afc03b589006368a9002da0014903b589006371a90203b5090012092a99a27602758335090003368900946e829619c1054511a00145e6704674a6740679e669466aa66a066b09618280907588711c6e9755ffff938575a12d468287907588711c6e9755ffff938505a139468287411106e497000000e78080010000411106e497000000e780a0000000411106e497b0ffffe780c0170000757106e5014730012948bd4821a89306f6ff13d547009a92a30f56fe0507368663fcf800aa879372f50013030003e3e002ff13037005e1bf13050008198d130610086370c5021755ffff9307a59e09462e85be8597000000e7800082aa60496182809305000897000000e78040660000757106e522e1a6fccaf8cef4d2f0d6ecdae8dee4e2e066fc6af86ef432892e8a014c814c81499715010003bb45d09715010083bb45d09715010083b445d000690c612ef008652aec13058a002ae01755ffff1305c5952ae8294d22e40da03305b6000345f5ff5915133515002300a4006265146d02758296ee8c6311051213f5f90f631b051063758901e9a8636c890d33058941b3058a014146637fc50063022c0d81463386d50003460600630da6098506e319d5fe75a013867500937686ff3386b640ad8e93b6160013371600d98ea1c20146930605ff02676297b387c5009c6313c4f7ffa58fda9733747401e18f8defb307c7009c6313c4f7ffa58fda9733747401e18f95e34106e3f9c6fc31a83387d500034707006307a7038506e319d6fe930605ffe3f9c6fa6304c5062264b386c50083c606006386a6010506e319c5fe05a0b286e296138c1600e3f026f5d29603c50600e31ba5f38149e28de28a39a04a8c8549e68dca8a63872c030345040001c96265146d11460275c265829611ed33869a41b3059a01e39a9aed0145f1bd4a8c2264f9b7014511a00545aa600a64e6744679a679067ae66a466ba66b066ce27c427da27d49618280411106e41b8605009306000802c26376d6002302b100054671a01bd6b50019ee13d665001366060c2302c10093f5f50393850508a302b1000946ada01bd6050115e613d6c5001366060e2302c10013964503699213060608a302c10093f5f503938505082303b1000d462da81396b50275921306060f2302c1001396e502699213060608a302c100139645036992130606082303c10093f5f50393850508a303b10011464c0097000000e780e0d9a26041018280397106fc907594712ae032f836f4886d906994658c612af032ec36e82ee41745ffff9305c57f0a85300097000000e780a0b2e27021618280086117030000670063d5411106e408611b8605009306000802c26376d6002302b100054671a01bd6b50019ee13d665001366060c2302c10093f5f50393850508a302b1000946ada01bd6050115e613d6c5001366060e2302c10013964503699213060608a302c10093f5f503938505082303b1000d462da81396b50275921306060f2302c1001396e502699213060608a302c100139645036992130606082303c10093f5f50393850508a303b10011464c0097000000e78060caa26041018280397106fc90759471986d32f836f43af0906994658c61086132ec36e82ee42ae01745ffff930525700a85300097000000e78000a3e27021618280357106ed22e926e54ae1cefcd2f8d6f42a840345050109c5833a04008544d5a0b2892e89033a840003654a03833a04009375450091e93336500163880a021745ffff9305855d35a063960a0483358a0203350a02946d9745ffff9385255c094682961dc5814a854469a81745ffff9305055b83368a0203350a02946e05068296854441e103b689014a85d28502968da803254a038544a303910283350a0203368a022ee432e8930571022eec83250a0303068a0383360a0003378a0083370a0103388a01aaceaecc2300c10636f43af83efcc2e02800aae403b689011745ffff1305c54faae82c104a85029619e9c6652665946d9745ffff9385055209468296aa8423089400850a233054012285ea604a64aa640a69e679467aa67a0d618280357106ed22e926e54ae1cefcd2f8d6f42a8403458500854a854419cd23049400a30454012285ea604a64aa640a69e679467aa67a0d6182803289ae89033a040003654a03834594001376450005e691cd83358a0203350a02946d9745ffff9385c54909468296854455f94e85d2850299aa846db785e183358a0203350a02946d9745ffff9385c54705468544829659f503254a038544a303910283350a0203368a022ee432e8930571022eec83250a0303068a0383360a0003378a0083370a0103388a01aaceaecc2300c10636f43af83efcc2e02800aae41745ffff1305053eaae82c104e85029915f9c6652665946d9745ffff9385454009468296aa8439bf397106fc22f826f44af02a841c7508719c6f3a89b684829722e8230ca10002e4a30c01002800a6854a8697000000e78060db22658345810139c50544b9e5834591017d1513351500c264b335b0006d8d05c103c54403118901ed8c748870946d9745ffff9385b53905460544829611ed8c748870946d9745ffff93856532054682962a8419a03334b0002285e2704274a274027921618280411106e497000000e78040920000757106e5014730012948bd4831a89306f6ff9377f50f13d547009a92a30f56fe0507368663fbf8001373f50093020003e36f03fd93027003d9bf13050008198d130610086370c5021745ffff9307053109462e85be8597f0ffffe7806014aa60496182809305000897000000e780a0f80000757106e5014730012948bd4831a89306f6ff9377f50f13d547009a92a30f56fe0507368663fbf8001373f50093020003e36f03fd93027005d9bf13050008198d130610086370c5021745ffff9307e52909462e85be8597f0ffffe780400daa60496182809305000897000000e78080f100001745ffff9306e53609462e85b68517f3ffff6700432e397106fc22f826f42e848c752ae40870946d9745ffff9385e5364546829622ec2300a10202e8a30001021745ffff1306653308082c0097000000e780a0c042658345010239c50544b9e5834511027d1513351500e264b335b0006d8d05c103c54403118901ed8c748870946d9745ffff9385f51e05460544829611ed8c748870946d9745ffff9385a517054682962a8419a03334b0002285e2704274a27421618280757106e5014730012948bd4821a89306f6ff13d547009a92a30f56fe0507368663fcf800aa879372f50013030003e3e002ff13037003e1bf13050008198d130610086370c5021745ffff9307651709462e85be8597f0ffffe780c0faaa60496182809305000897000000e78000df0000797106f422f026ec4ae84ee42a8404690865ae893309b640058d6363250308602695ce854a8697f00000e78060dfca9404e8a2700274e2644269a269456182802285a6854a8697000000e780c0000468f9b75d7186e4a2e026fc2e966368b6042a8408659314150063639600b284a14563e39500a14493c5f4fffd9119c5106032f0054632f42af811a002f428001410268697000000e780e003a265426581cdfd55fe158505630ab50009ed97b0ffffe780408a000008e004e4a6600664e27461618280626597b0ffffe78000880000011106ec22e826e44ae03289aa8499cd2e84886605c18c6a91cd88624a8697b0ffffe780808405e180e419a023b40400854521a8630409024a85a28597b0ffffe780a08175d1814588e423b824018ce0e2604264a264026905618280228565f5e1b703e6450308619376060191ea1376060209ee0345050017f3ffff670063d00305050017030000670023d10305050017030000670043c903e6450308619376060189ea1376060219ea086117f3ffff670023cd086117f3ffff67006359086117030000670003e0411106e422e02a8411c96347040289c9228597a0ffffe780407909a8054501a88545228597a0ffffe780a07619c9a285a26002644101828097a0ffffe78000780000228597a0ffffe780a07600005d7186e4a2e026fc4af84ef452f0ae898c750461006903b50902946d9745ffff938525f00546054982964ee42308a100a308010005c417050000930965f1138a140026ec28002c084e8697000000e780e0a17d14d28465f40345010101ed22650c750871946d9745ffff9385f5ef054682962a894a85a6600664e2744279a279027a61618280797106f422f026ec4ae84ee42a8904690865058d2e84636fb50283390900894533859900636cb4007d148145228697f00000e78040aba2943385990023000500850423389900a2700274e2644269a269456182804a85a685228697000000e780e0008334090155bf5d7186e4a2e026fc2e966368b6042a8408659314150063639600b284a14563e39500a14493c5f4fffd9119c5106032f0054632f42af811a002f428001410268697000000e780e003a265426581cdfd55fe158505630ab50009ed97a0ffffe7802062000008e004e4a6600664e27461618280626597a0ffffe780e05f0000011106ec22e826e43284aa8499cd88660dc18c6a99cd8862228697a0ffffe780a05c19ed85458ce431a823b40400854511a88545228597a0ffffe780e0597dd1814588e480e88ce0e2604264a26405618280411106e422e02a8408617d1508e005e90c70086c8c6182950870086511c5086c97a0ffffe780a056087811c5087497a0ffffe780c05508647d1508e409c5a2600264410182802285a2600264410117a3ffff6700c3535d7186e4a2e026fc4af84ef452f056ec83ba0501368a3289aa8963e3da00d28a806108687de1286c7d5610e8637c55010870106c98651c6d4e85b2854a86d286829761a08465306463edc400b386540163ee96082c683307b600636ec7086376d70208700c6c1074147c1c6d0a85268782970345010069e9a26563e8550f286c2ce824e426866367b50eb3b6c400918c33359500558d49e5338554016363950463e7a5080c7c63eca508b3059540639745090c74a6954a85528697f00000e780809623b45901238009000868050508e8a6600664e2744279a279027ae26a616182801745ffff130525e411a81745ffff130585e329a01745ffff1305e5e2f14597f0ffffe780800400001745ffff1305b5d89745ffff9386a5d9c1450a8689a01745ffff1305a5e69305f002d1bf1745ffff1305b5e893052003d9b7528597000000e780e08a00001745ffff1305a5039745ffff938645db9305b0021306710197f0ffffe780801900001745ffff130565dd71b71745ffff130585de9305e00241b7034505000e051746ffff1306c6362a969746ffff9386263b369598751062146188711c6fb6858287411110650c69b29563edc50008611069fd568582637dd60028616369b502410182801745ffff130505aba14535a01745ffff130545cf9745ffff938645d0e145300097f0ffffe780c01000001745ffff130555df9305600297f0ffffe78060f40000797106f422f0aa8502c2280050009146114497000000e78020de0345810011e942656319850203654100a2700274456182801745ffff130545f49745ffff9386e5cb9305b0021306f10197f0ffffe780200a00001745ffff130515dbb54597f0ffffe780e0ed0000411106e497000000e78040f98d4563f7a50009817d15a260410182801745ffff1305e5d8b94597f0ffffe780e0ea0000197186fca2f8a6f4caf0ceecd2e8d6e4dae05efc03bb050003370b00806594692a89130517002330ab0065c95ae409072330eb007dc3b28a36f85af02e8597000000e780a0f29305440063ea850caa892ef4081097000000e780c0f763ffaa02aa84938b1a0013952b002295636e850a2af4081097000000e78040ef2a8a63999b02330544016366850a2ae863f649051745ffff130525ddc1a015452304a900233009005a8597000000e78000c6b1a08a0a33858a002105636285082af4081097000000e78080eab305440163ed8506aa892ee8636e4507338549412aec280097000000e78060e26265c26522662338a9002334b9002330c9005a8597000000e780a0c0e6704674a6740679e669466aa66a066be27b09618280000000001745ffff130545d40da81745ffff1305a5d325a01745ffff130505d339a81745ffff130565d211a81745ffff1305c5d129a01745ffff130525d19305b00297f0ffffe78080d40000797106f422f0906118629465050718e20dcf2a841385460032e4636ad5022ae82e8597000000e78000de2aec280097000000e78020d76265c265226608e80ce410e0a270027445618280000000001745ffff1305e5ca9305b00297f0ffffe78040ce0000397106fc22f826f42a8402e408083000a146a144a28597000000e780c0b70345010105e16265631f9502a264086097000000e780e0b02685e2704274a274216182801745ffff130525cd9745ffff9386c5a49305b0021306710297f0ffffe78000e300001745ffff1305a5b5b94597f0ffffe780c0c60000397106fc22f826f42a84a307010008081306f10085468544a28597000000e78000b0034501010de16265631095048304f100086097000000e78000a92685e2704274a274216182801745ffff130545c59745ffff9386e59c9305b0021306710297f0ffffe78020db00001745ffff130585afb54597f0ffffe780e0be00005d7186e4a2e026fc4af8ae842a898c69054632e002e402e889c90a8597000000e780208f0266426411a001442808a685a28697000000e780a0a6034581011de5027563168504c2652266826688602338b9002334c9002330d900a6600664e27442796161170300006700239e1745ffff130525bb9745ffff9386c5929305b0021306f10297f0ffffe78000d100001745ffff130535a6c94597f0ffffe780c0b40000011106ec22e826e49c692a84637df700b384e74063e3d400b684b306970063ede60263f7d7001545a300a400054531a8998e639dd4028c61ba953285268697e00000e780e03d014504e42300a400e2604264a264056182801745ffff1305658cf14597f0ffffe78000ae00002685b68597f0ffffe780603700005d7186e4a2e026fc4af84ef452f02e8483b905012a896145a14597a0ffffe78020e959c1aa84086888e8086488e4086088e0054a52e402e802ec1314ba002800a28597f0ffffe780007b13050006a14597a0ffffe780c0e531c923304501233445012338050004ed9745ffff938545980cf1a2650cf5c2650cf9e2650cfd23303505233405042338050420ed23340900233839012330a900a6600664e2744279a279027a61618280614519a01305000697a0ffffe780c0e100000c6591c5086117a3ffff670043df8280397106fc22f826f44af09376f60f1307f00f2a89638fe6041b04160002ec02e802e402e0131584036d9113060002098e8a84aa94aa95268597e00000e780002a1375740009c9838504007d563315a6006d8d2380a4008a85130600024a8597e00000e780a027e2704274a274027921618280130600024a858145e2704274a2740279216117e30000670063182a860345050283c605023337d500358d3335a000b306e040558d0de5fd057d06815695c20345060003c70500b337e500398d3335a0003307f040598dfd157d16850665d18280014582805d7186e4a2e026fc4af8ae84806590612a892800a28597e0ffffe78080b30345810019c5426529e109452300a90029a805040dc09305910080e4130610024a8597e00000e780201ca6600664e2744279616182801745ffff1305058cf14597f0ffffe780a08c000097f0ffffe780c0a80000306115ce14610c653337d00093b715007d8f7d1630e115c7106d0c699306050109c683b505227d166dfe0146014723b4060023b00600854614e10ce531a08145b1a8b5ca1869106d83d6a5216374d600ae8621a883b60521a1c603d6852183d7a6210507b685e377f6fe1308160001cf0e083698833708227d1701c783b70722e5bf014811a0b68793050003b305b602b6951ce523380500233c05012e8582801735ffff1305457d9305b00297f0ffffe780a08000001735ffff1305e57bedb7411106e413050022c14597a0ffffe78000bd01c5a260410182801305002297a0ffffe780c0bd0000411106e413050028c14597a0ffffe78080ba01c5a260410182801305002897a0ffffe78040bb00001d7186eca2e8a6e4cae04efc52f856f45af05eec62e866e46ae03e893a8ab689b28aae8b2a84035ca52193841500139b55002a9b139d4500b30cbc40637b9c00130600025a85d68597e00000e780800381a013955400229513965c00da8597e00000e7800047130600025a85d68597e00000e780200113050416b305a50113964400329513964c0097e00000e7806044930a1c00229d23344d1723303d1793092c00130a042213852b00139b3400637c3501b3056a010e05529513963c0097e00000e78000415a9a23302a01231d542163f434038e0ba29b13858b22b305804109461461239c9620850423b88620b38695002105e397c6fee6604664a6640669e279427aa27a027be26b426ca26c026d256182800358a5212e86814593125800aa929303f5011303f601054e63055504938815001305050201579a869e8715cf83ce060003c6070033bfce0033c6ce00b33ec0003306e0413366d601fd17fd16050771de1376f60f631ac60193830302c685e31f55fac28511a0014e72858280457186e7a2e326ff4afb4ef752f356ef5aeb5ee762e3e6feeafaeef62e8a83bb050083b90501b28a2a8b03d9ab21139559005e9583459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18d2ef483451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2ef083459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2eec83451500034605008346250003473500a205d18dc2066207d98ed58d034655008346450003476500834775002206558e4207e2075d8f598e0216d18d2ee8938c190093955c00de9513c6f9ff330426011316540097e00000e780c02093850b16139549002e950465033c050013964c00b2951316440097e00000e780a01e7d3913150903239d2b21033a8a0041919545637bb51a2819de8552869760ffffe780a0736a7556e026e405cd85456317b5068001080113068003a28597e00000e78080d56a65aa750355a52183d5a5212e950505b1456376b50408180c01014605a88001a80013068003a28597e00000e78080d20675c6750355a52183d5a5212e950505b1456372b5040818ac000546ce8697000000e780604899a80e65ae650da0081a13068003a28597e00000e780a0ce081a854597000000e780c0153665d6652af82efccee025a0081a13068003a28597e00000e78020cc081a854597000000e7802072766596752af82efce6e0c27b627a03b60b21866971c613041a00930a010c914c314d954d05498354a62163eb9c0a2819b28522869760ffffe780c0636a751dcd631b2509a81913068003d68597e00000e78020c6526592750355a52183d5a5212e950505636ea503b3859d40a81997000000e780e00b01465df69da0a81913068003d68597e00000e780a0c2526592750355a52183d5a5212e9505056373a503081a13068003d68597e00000e78060c0081a97100000e78080932a862e8425f605a0b3859d40a81997000000e7802065014631fa31a089e4054582652380a500a264227582756266c266233cab002338bb002334cb002330db0023308b0323349b0223387b03233c4b0323303b05be601e64fa745a79ba791a7afa6a5a6bba6b1a6cf67c567db67d79618280317106fd22f926f54af14eed52e956e55ae1defce2f8e6f4eaf0eeec6383052a2e892a8a833b850183d5ab21338425012d45636e85282ef4033b8a020355ab21636e252933052541239d8b202ae4231dab20930af9ff93945a0093090b1613954a002ae84e9583350a01833d0a00106532f008612aec139555006e959205ae9d83459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18daee483451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18daee083459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2efc83451500034605008346250003473500a205d18dc206620703465500d98ecd8e83454500220603476500834775004d8e268cb3059b004207e2075d8f598e0216558e32f81306000297e00000e780e0e403bd0d1683bc8d16626523b0ad16027523b4ad16a28da274139554005e950c181306000297e00000e780409d13840b16139544002295233495018504b3859d402330a501639cba10139554005e95da85628697e00000e780609a139544002295ce85426697e00000e780409993155900da95226c13165c005a8597e00000e780c0dc93154900ce9513164c004e8597e00000e78080db83350a0203350a03adcd79c113040b22139534005e951305052293193900a2854e8697e00000e7800094b305340113163c002106228597e00000e780a0d7a27c63f0bc038e0cde9c13858c220c61239c9520850423b875217d192105e31809fe7d556301ac020145050c0c601306150023b86521239ca52021043285e317ccfe11a039e5ea704a74aa740a79ea694a6aaa6a0a6be67b467ca67c067de66d296182801735ffff13050516ed4505a81735ffff1305151f930520030da01735ffff1305552111a81735ffff1305f50d29a01735ffff1305751a9305800297e0ffffe780c0fa0000317106fd22f926f54af14eed52e956e55ae1defce2f8e6f4eaf0eeec806d035da4216a8701c698750357a721636cd72832f036f42af883ba850203dcaa21930b1d0033868b012d456365c528846188652ae803b9050188712aec03dba42132e4231dc42013155900269583459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18daee883451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18daee483459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18daee083451500034605008346250003473500a205d18dc2066207d98ed58d034655008346450003476500834775002206558e4207e2075d8f598e0216d18d2efc930d190093955d00a6959349f9ffda991396590097e00000e78040b513155d0022952c181306000297d00000e780206f13955b00229513165c00d68597d00000e780e06d93850416131549002e95033a0500833c850013964d00b2951396490097e00000e78080b01305041693154d00aa9523b4950123b0450193850a1613964b00329513164c0097d00000e78020699385042213953d002e950e09ca95c1051396390097e00000e78040ac63f06d032699130589220c6113861d0023b89520239cb5212105b28de317cbfe0395a4217d358545239da420426563f3a50413953b0022951305052293850a2213163c00210697d00000e780806222656372ad02050c0e0d229d13058d22de851061231cb6208505233886207d1c2105e3180cfe02759334150056859790ffffe7804010fd1433f57401a2752e95c27580e1626690e588e9ea704a74aa740a79ea694a6aaa6a0a6be67b467ca67c067de66d296182801735ffff1305f5f49305100939a01735ffff130525fd9305a00297e0ffffe78040cc0000717106f522f126ed4ae94ee552e1d6fcdaf8def4e2f0e6eceae8eee4638605262e8b2a890075835ca421e6952d456363b526033c89018354ac2163e46427338d6441231dac212ee4231db42013155b00229513965c00a28597e00000e780a0989309041613154b004e9513964c00ce8597e00000e7802097930b1d00b38a74411305fbff6396aa2293955b00e295139a5a002285528697d00000e780e04f93040c1693954b00a695920a4e85568697d00000e780604e13154d00269583350901833d0900106532ec08612ae8139555006e959205ae9d83459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18d2efc83451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2ef883459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2ef483451500034605008346250003473500a205d18dc20662070346550083474500d98ecd8e22065d8e034765008347750093155d00e2954207e2075d8f598e0216558e32f01306000297e00000e780a08003bd0d1683b48d16426523b0ad16626523b4ad16330544010c101306000297d00000e7806039d69923b4990023b0a9018335090203350903a1c945c1930404220e0b3385640113963c002106a68597d00000e780407b8e0be29b93850b2226855a8697d00000e780203581452265050590609386150023388620231cb620a104b685e317d5fe11a029e9aa700a74ea644a69aa690a6ae67a467ba67b067ce66c466da66d4d6182801735ffff1305c5baed4515a81735ffff1305b5bb930530031da01735ffff130505be9305700221a81735ffff130575b229a01735ffff1305f5be9305800297e0ffffe780409f0000357106ed22e926e54ae1cefcd2f8d6f4daf0deece2e8e6e4eae06efc033a850183398502835aaa2103dba92113841a0033066401ad4563e1c526033d0500833c050108652ae8035cad2132e4231dca2013955c006a9583459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18d2ef883451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2ef483459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2ef083451500034605008346250003473500a205d18dc2066207d98ed58d034655008346450003476500834775002206558e4207e2075d8f598e0216d18d2eec93841c0093955400ea9593cdfcffe29d13965d0097d00000e780005b13955a0052952c081306000297d00000e780e01413155400529513165b00ce8597d00000e780a01393050d1613954c002e9503390500833b850013964400b29513964d0097d00000e780405613050a1693954a00aa9523b4750123b025019385091613164400329513164b0097d00000e780e00e93050d22139534002e958e0ce695c10513963d0097d00000e780005263f08403ea9c13858c220c611386140023b8a521239c95202105b284e317ccfe0315ad217d358545231dad20c26463f29504131534005295130505229385092213163b00210697d00000e7804008226563f1aa02050b8e0ad29a13858a220c61239c8520050423b845217d1b2105e3180bfe4e859790ffffe78080b66a85a685ea604a64aa640a69e679467aa67a067be66b466ca66c066de27d0d6182801735ffff130545a59305a00297d0ffffe78060740000411106e413058072a1459790ffffe78060b101c5a26041018280130580729790ffffe78020b20000411106e413058078a1459790ffffe780e0ae01c5a26041018280130580789790ffffe780a0af00001d7186eca2e8a6e4cae04efc52f856f45af05eec62e866e43a89b689328a2e8b2a84835b655b1305855b938415009605da95b30ab500338c6b4163fb9b00130610025685d28597d00000e78000f8a9a09395540026952e9513165c006296d68597d00000e780403b130610025685d28597d00000e78060f51305840013064008b305cb02aa95b386c40236953306cc0297d00000e7804038138a1b00130540083305ab022295210513064008ce8597d00000e78080f193892b00930a847213052b00939c3400637c3501b3859a010e05569513163c0097d00000e780e033e69a23b02a01231b445b63f334030e0b229b13050b73b305704109461461239a965a850480e2b38695002105e398c6fee6604664a6640669e279427aa27a027be26b426ca26c25618280397106fc22f826f44af04eec52e856e48359655b2e8a9305855b93945900ce947d54054995c4938a1502528597f0ffffe78060c29384f4fd1375f50f0504d685e30225ff9305f00f6305b500014911a04e844a85a285e2704274a2740279e269426aa26a21618280130101ce233c1130233881302334913023302131233c312f2338412f2334512f2330612f233c712d2338812d2334912d2330a12d233cb12b2e8c83bb050003bb05013289aa8903da6b5b13848b5b13155b005a95b30ca400a80b13061002e68597d00000e78060dd930a1b0093955a005694a2951345fbffb3044501139654002696668597d00000e7800020930c400833059b033384ab00130d84001305911f13064008ea8597d00000e78000d99305c408338694036a8597d00000e780c01c1b05faff239bab5a033a8c004215135405032811ac0b1306500a97d00000e780c0d50a852c111306500a97d00000e780c0d41545637da41a2811de85528697000000e78060202a7505cd85456317b5060019081313068003a28597d00000e780c0d17a75be650355655b83d5655b2e950505b1456376b504880a0c13014605a80019a81213068003a28597d00000e780c0ce1a65da650355655b83d5655b2e950505b1456372b504880aac120546da8697000000e780004ca9a84a75ea750da0a80b13068003a28597d00000e780e0caa80b854597000000e780601d5e75fe75aaeaaeeedaf235a0a80b13068003a28597d00000e78060c8a80b854597000000e780a06b0335012083358120aaeaaeeed6f2d66b766a03b60b00167b69ca93041a00930a010b914d314c954c054d0354665b63ee8d0a2811b285268697000000e78080102a7529c1631fa509080513068003d68597d00000e78020c2033581298335812a0355655b83d5655b2e95050563608505b3858c40080597000000e780001301464df6a5a0080513068003d68597d00000e78060be033581298335812a0355655b83d5655b2e95050563738503a80b13068003d68597d00000e780e0bba80b97100000e78020882a86ae8425f239a8b3858c40080597000000e780e05d014631f629a001e405452300a9008a851306500a4e8597d00000e78000b823b4790b23b8490b23bc690b833081310334013183348130033901308339812f033a012f833a812e033b012e833b812d033c012d833c812c033d012c833d812b13010132828094619dc683d7455b130816009dc71387f7ff93173700b69783b787722330050014e52338050118ed1cf110f50cf92da00ce510e989450ce1828003d7665b19cf03b7067385471ce114e523380501233c05000cf110f518f910fd828097d0ffffe780803c0000130101d92334112623308126233c9124233821252334312523304125233c5123233861232334712323308123233c91212338a1212334b121638505242e89aa8b033d850103546d5bb304b4002d456360952422ec83bc8b0203d56c5b63602525330a2541231b9d5a239b4c5b930df9ff93898c5b13955d006e952ae4338ba900938a8c0013044008b3858d022ee8d69528101306400897d00000e78060a303b50b0183b50b0013165500b386a500369626f09304865b330585022e95130c8500081913061002a68597d00000e78040a0130610022685da8597d00000e78020e49304110d130640082685e28597d00000e780009e2c1013064008628597d00000e780009da80a0c191306100297d00000e780009c080313064008a68597d00000e780009b130b8d5b626c13155c00b3058b012e95ac0a1306100297d00000e780209993048d0033058c0226950c031306400897d00000e780a09713041c000275018d6392ad1413155400229b5a95ce85226697d00000e780a095130b4008330564032695d685426697d00000e7804094131559004a95b385a90013165a0052964e8597d00000e78080d7b3056903d69533066a03568597d00000e78040d683b50b0203b50b03c1c165c5d28a93848c72131534006a951305857293193900a6854e8697d00000e780a08eb385340113163a002106268597d00000e78040d202756371ac02131a3c006a9a13050a730c61239a855a050423b0a5017d192105e31809fe7d556382aa02814513851a0090609386150023309601231ab65aa104b685e317d5fe11a02de58330812603340126833481250339012583398124033a0124833a8123033b0123833b8122033c0122833c8121033d0121833d81201301012782801725ffff1305a50eed4505a81725ffff1305b517930520030da01725ffff1305f51911a81725ffff1305950629a01725ffff130515139305800297d0ffffe78060f30000697106f622f226ee4aea4ee652e2d6fddaf9def5e2f1e6edeae9eee583bd850103dc6d5b628701c698750357675b636ad71e32f036f42af883ba850283dc6a5b130b1c0033069b012d456363c51e846188652ae888712aec83b9050183db645b32e4239bcd5a1384845b139559004e95330da400880013061002ea8597c00000e780a07813891900931559004a94a29513caf9ff5e9a52fc13165a0052966a8597d00000e78040bb13848d5b13155c00b30584012e958c001306100297c00000e780a07493858a5b13155b005a94229513965c00669697c00000e7800073130d40083385a9033384a400628a5a8c668bd68c930a8400880013064008d68597c00000e78080709305c40862753306a5035685e68ada8c628b97d00000e780c0b313848d003305aa0322958c001306400897c00000e780606d93858a003305ac0322953386ac0397c00000e780006c93858472131539002e958e09ce95c10562760e0697d00000e78020af637f7901a699138509730c611306190084e1239a255b21053289e398cbfe0395645b7d358545239ba45a426563f4a50413153b006e951305857293858a7213963c00210697c00000e780806522656373aa02850c131c3a006e9c13050c73da851061231ab65a85052330b601fd1c2105e3980cfe02751334150056859780ffffe78020137d1433756401a2752e95c27523b0b501626690e588e9b2701274f2645269b269126aee7a4e7bae7b0e7cee6c4e6dae6d556182801725ffff1305b5f79305100939a01725ffff1305e5ff9305a00297d0ffffe78000cf0000130101d92334112623308126233c9124233821252334312523304125233c5123233861232334712323308123233c91212338a1212334b121638705202e8caa8b0075035d645bea952d456364b52003bb8b01835a6b5b63e58a21338a8a41231b4b5b2ee8231bb45a1309845b13155c0062954a9513165d006a96ca8597d00000e780209993098400930c400833059c034e9533069d03ce8597d00000e7806097930d1a00b384ba411305fcff6391a41cda8a130b8b5b93955d003305bb01aa95139554003306950032f04a8597c00000e780404f56e4a10ab3859d03d6953386940332ec4e8597c00000e780a04d13155a00529b2a9bb3059a03d69528101306400897c00000e780e04b03b50b0183b50b0013165500b386a50036969304865b330595032e95930c8500081913061002a68597c00000e780e048130610022685da8597d00000e780c08c9304110d130640082685e68597c00000e780a0462c1013064008668597c00000e780a045a80a0c191306100297c00000e780a044080313064008a68597c00000e780a04302754a95ac0a1306100297c00000e780804262654e950c031306400897c00000e780604183b50b0203b50b03a1c955cd930484720e0c3385840113163d002106a68597d00000e780e0838e0d2265aa9d93858d722685628697c00000e780a03d81454265050590609386150000e2231ab65aa104b685e318d5fe11a03de58330812603340126833481250339012583398124033a0124833a8123033b0123833b8122033c0122833c8121033d0121833d81201301012782801725ffff1305a5c1ed4515a81725ffff130595c2930530031da01725ffff1305e5c49305700221a81725ffff130555b929a01725ffff1305d5c59305800297d0ffffe78020a600006d7106e622e2a6fdcaf9cef5d2f1d6eddae9dee5e2e166fd6af96ef5033a850183398502035b6a5b83db695b13041b0033067401ad4563ebc51a833c05000c652eec833d050103dd6c5b32e0231bca5a13898c5b13955d006e95b30aa900081013061002d68597c00000e780c02c93841d00939554002699ca9513c9fdff6a99131659004a96568597c00000e780806f930a8a5b13155b00b3856a012e950c101306100297c00000e780e0289385895b13155400a29a569513965b005e9697c00000e7804027130c400833858d03b38aac005ee4ce8b93898a00081013064008ce8597c00000e78000259385ca08330689034e8597c00000e780c06893098a005ae833058b034e950c101306400897c00000e7804022de8a93858b00a26b330584034e9533868b0397c00000e780a02093858c72139534002e958e0dee95c1051316390097c00000e780c06363f0a403e69d13850d730c611386140023b09501239a955a2105b284e317cdfe03956c5b7d358545239bac5ae264426b63f295041315340052951305857293858a7213963b00210697c00000e780e01902656371ab02850b0e0b529b13050b730c61239a855a050423b04501fd1b2105e3980bfe56859780ffffe78020c86685a685b2601264ee744e79ae790e7aee6a4e6bae6b0e6cea7c4a7daa7d516182801725ffff1305e5b69305a00297d0ffffe78000860000130101dc233c1122233881222334912223302123233c3121233841212334512123306121deffe2fbe6f7eaf3eeefd54bae8a63f575052a8c094563e9aa0005466285d68597300000e78060e98330812303340123833481220339012283398121033a0121833a8120033b0120fe7b5e7cbe7c1e7dfe6d130101248280b68cb2892afc930d7113054d0545aae856f8627c1b850c0019e16f20f00613751d0019e16f10b07d466813db2a0013171b00b308670113051003637955231303fbff93021b0013166b00629603459601834586018346a6018347b60122054d8dc206e207dd8e558d8345d6018346c6018347e6018344f601a205d58dc207e204c58fdd8d82154d8d2af90345160183450601834626018347360122054d8dc206e207dd8e558d83455601834646018347660183447601a205d58dc207e204c58fdd8d82154d8d2af503459600834586008346a6008347b60022054d8dc206e2078345d6008344c600dd8e558da205cd8c8346e6008347f60093156300e295c206e207dd8ec58e8216558d2af1034516008346060083472600834436002205558dc207e204c58f5d8d83465600834746008344660003467600a206dd8ec2046206458e558e0216518d2aed03c5950103c6850183c6a50183c7b5012205518dc206e207dd8e558d03c6d50183c6c50183c7e50183c4f5012206558ec207e204c58f5d8e0216518d2afa03c5150103c6050183c6250183c735012205518dc206e207dd8e558d03c6550183c6450183c7650183c475012206558ec207e204c58f5d8e0216518d2af603c5950003c6850083c6a50083c7b5002205518dc206e207dd8e558d03c6d50083c6c50083c7e50083c4f5002206558ec207e204c58f5d8e0216518d2af203c5150003c6050083c6250083c735002205518dc206e207dd8e558d03c6550083c6450083c7650083c575002206558ec207e205dd8dd18d82154d8d2aee01559305710b6e8605c583c60500834706007d16fd150505e388f6feb3b3f60063f9f6009a875a8331a081436f10c0168143da8713956200629503469501834685018344a5010344b5012206558ec2046204458c418e8346d5018344c5010344e5018345f501a206c58e4204e205c18dd58d8215d18d2ef983451501034605018346250183443501a205d18dc206e204c58ed58d034655018346450183446501034475012206558ec2046204458c418e0216d18d2ef583459500034685008346a5008344b500a205d18dc206e2040346d5000344c500c58ed58d2206518c8346e5008344f500139667006296c206e204c58ec18e8216d58d2ef183451500834605008344250003443500a205d58dc2046204458cc18d83465500834445000344650003457500a206c58e42046205418d558d02154d8d2aed03459601834586018346a6018344b60122054d8dc206e204c58e558d8345d6018346c6018344e6010344f601a205d58dc2046204458cc18d82154d8d2afa0345160183450601834626018344360122054d8dc206e204c58e558d83455601834646018344660103447601a205d58dc2046204458cc18d82154d8d2af603459600834586008346a6008344b60022054d8dc206e204c58e558d8345d6008346c6008344e6000344f600a205d58dc2046204458cc18d82154d8d2af20345160083450600834626008344360022054d8dc206e204c58e558d83455600834646008344660003467600a205d58dc2046206458ed18d82154d8d2aee01551306710b130471130dc183440600834604007d147d160505e388d4fe63e3d400be8233b5d400aa93968713956700629583459501034685018346a5018344b501a205d18dc206e204c58ed58d0346d5018346c5018344e5010344f5012206558ec2046204458c418e0216d18d2ef983451501034605018346250183443501a205d18dc206e204c58ed58d034655018346450183446501034475012206558ec2046204458c418e0216d18d2ef583459500034685008346a5008344b500a205d18dc206e2040346d5000344c500c58ed58d2206518c8346e5008344f500131663006296c206e204c58ec18e8216d58d2ef183451500834605008344250003443500a205d58dc2046204458cc18d83465500834445000344650003457500a206c58e42046205418d558d02154d8d2aed03459601834586018346a6018344b60122054d8dc206e204c58e558d8345d6018346c6018344e6010344f601a205d58dc2046204458cc18d82154d8d2afa0345160183450601834626018344360122054d8dc206e204c58e558d83455601834646018344660103447601a205d58dc2046204458cc18d82154d8d2af603459600834586008346a6008344b60022054d8dc206e204c58e558d8345d6008346c6008344e6000344f600a205d58dc2046204458cc18d82154d8d2af20345160083450600834626008344360022054d8dc206e204c58e558d83455600834646008344660003467600a205d58dc2046206458ed18d82154d8d2aee01551306710b9304711315c10344060083c60400fd147d160505e308d4fe6363d4003e833335d400aa931a8b11a03e8b9304f7ff9362170013156700629583459501034685018346a5018347b501a205d18dc206e207dd8ed58d0346d5018346c5018347e5010344f5012206558ec2076204c18f5d8e0216d18d2ef983451501034605018346250183473501a205d18dc206e207dd8ed58d034655018346450183476501034475012206558ec2076204c18f5d8e0216d18d2ef583459500034685008346a5008347b500a205d18dc206e2070346d5000344c500dd8ed58d2206518c8346e5008347f500139664006296c206e207dd8ec18e8216d58d2ef183451500834605008347250003443500a205d58dc2076204c18fdd8d83465500834745000344650003457500a206dd8e42046205418d558d02154d8d2aed03459601834586018346a6018347b60122054d8dc206e207dd8e558d8345d6018346c6018347e6010344f601a205d58dc2076204c18fdd8d82154d8d2afa0345160183450601834626018347360122054d8dc206e207dd8e558d83455601834646018347660103447601a205d58dc2076204c18fdd8d82154d8d2af603459600834586008346a6008347b60022054d8dc206e207dd8e558d8345d6008346c6008347e6000344f600a205d58dc2076204c18fdd8d82154d8d2af20345160083450600834626008347360022054d8dc206e207dd8e558d83455600834646008347660003467600a205d58dc20762065d8ed18d82154d8d2aee01551306710b9306711315c18347060003c40600fd167d160505e38887fe33b58700aa9363f58700a686ba8411a0ba8613956200629583459501034685010347a5018347b501a205d18d4207e2075d8fd98d0346d5010347c5018347e5010344f5012206598ec2076204c18f5d8e0216d18d2ef983451501034605010347250183473501a205d18d4207e2075d8fd98d034655010347450183476501034475012206598ec2076204c18f5d8e0216d18d2ef583459500034685000347a5008347b500a205d18d4207e2070346d5000344c5005d8fd98d2206518c0347e5008347f5001396660062964207e2075d8f418f0217d98d2ef183451500034705008347250003443500a205d98dc2076204c18fdd8d0347550083474500034465000345750022075d8f42046205418d598d02154d8d2aed03459601834586010347a6018347b60122054d8d4207e2075d8f598d8345d6010347c6018347e6010344f601a205d98dc2076204c18fdd8d82154d8d2afa0345160183450601034726018347360122054d8d4207e2075d8f598d83455601034746018347660103447601a205d98dc2076204c18fdd8d82154d8d2af603459600834586000347a6008347b60022054d8d4207e2075d8f598d8345d6000347c6008347e6000344f600a205d98dc2076204c18fdd8d82154d8d2af20345160083450600034726008347360022054d8d4207e2075d8f598d83455600034746008347660003467600a205d98dc20762065d8ed18d82154d8d2aee01551306710b130771130dc103440600834707007d177d160505e308f4fe6363f400b6823335f400aa93968613956600629583459501034685010347a5018347b501a205d18d4207e2075d8fd98d0346d5010347c5018347e5010344f5012206598ec2076204c18f5d8e0216d18d2ef983451501034605010347250183473501a205d18d4207e2075d8fd98d034655010347450183476501034475012206598ec2076204c18f5d8e0216d18d2ef583459500034685000347a5008347b500a205d18d4207e2070346d5000344c5005d8fd98d2206518c0347e5008347f5001396640062964207e2075d8f418f0217d98d2ef183451500034705008347250003443500a205d98dc2076204c18fdd8d0347550083474500034465000345750022075d8f42046205418d598d02154d8d2aed03459601834586010347a6018347b60122054d8d4207e2075d8f598d8345d6010347c6018347e6010344f601a205d98dc2076204c18fdd8d82154d8d2afa0345160183450601034726018347360122054d8d4207e2075d8f598d83455601034746018347660103447601a205d98dc2076204c18fdd8d82154d8d2af603459600834586000347a6008347b60022054d8d4207e2075d8f598d8345d6000347c6008347e6000344f600a205d98dc2076204c18fdd8d82154d8d2af20345160083450600034726008347360022054d8d4207e2075d8f598d83455600034746008347660003467600a205d98dc20762065d8ed18d82154d8d2aee01551306710b1307711315c183470600034407007d177d160505e38887fe63e38700b68433b58700aa93268711a036871383f8ff9382180013956800629583459501034685018346a5018347b501a205d18dc206e207dd8ed58d0346d5018346c5018347e5018344f5012206558ec207e204c58f5d8e0216d18d2ef983451501034605018346250183473501a205d18dc206e207dd8ed58d034655018346450183476501834475012206558ec207e204c58f5d8e0216d18d2ef583459500034685008346a5008347b500a205d18dc206e2070346d5008344c500dd8ed58d2206d18c8346e5008347f500131663006296c206e207dd8ec58e8216d58d2ef183451500834605008347250083443500a205d58dc207e204c58fdd8d83465500834745008344650003457500a206dd8ec2046205458d558d02154d8d2aed03459601834586018346a6018347b60122054d8dc206e207dd8e558d8345d6018346c6018347e6018344f601a205d58dc207e204c58fdd8d82154d8d2afa0345160183450601834626018347360122054d8dc206e207dd8e558d83455601834646018347660183447601a205d58dc207e204c58fdd8d82154d8d2af603459600834586008346a6008347b60022054d8dc206e207dd8e558d8345d6008346c6008347e6008344f600a205d58dc207e204c58fdd8d82154d8d2af20345160083450600834626008347360022054d8dc206e207dd8e558d83455600834646008347660003467600a205d58dc20762065d8ed18d82154d8d2aee01551306710b9304711315c18346060083c70400fd147d160505e388f6fe33b5f600aa9363f5f6001a86468311a0468613956200629583459501834685018347a5018344b501a205d58dc207e204c58fdd8d8346d5018347c5018344e5010344f501a206dd8ec2046204458cc18e8216d58d2ef983451501834605018347250183443501a205d58dc207e204c58fdd8d83465501834745018344650103447501a206dd8ec2046204458cc18e8216d58d2ef583459500834685008347a5008344b500a205d58dc207e2048346d5000344c500c58fdd8da206c18e8347e5000344f50093146600e294c2076204c18fdd8e8216d58d2ef183451500834605008347250003443500a205d58dc2076204c18fdd8d83465500834745000344650003457500a206dd8e42046205418d558d02154d8d2aed03c5940183c5840183c6a40183c7b40122054d8dc206e207dd8e558d83c5d40183c6c40183c7e40103c4f401a205d58dc2076204c18fdd8d82154d8d2afa03c5140183c5040183c6240183c7340122054d8dc206e207dd8e558d83c5540183c6440183c7640103c47401a205d58dc2076204c18fdd8d82154d8d2af603c5940083c5840083c6a40083c7b40022054d8dc206e207dd8e558d83c5d40083c6c40083c7e40003c4f400a205d58dc2076204c18fdd8d82154d8d2af203c5140083c5040083c6240083c7340022054d8dc206e207dd8e558d83c5540083c6440083c7640083c47400a205d58dc207e204c58fdd8d82154d8d2aee01559304710b130471130dc183c70400834604007d14fd140505e388d7fe63e3d700b28233b5d700aa93168613156600629583459501834685018347a5018344b501a205d58dc207e204c58fdd8d8346d5018347c5018344e5010344f501a206dd8ec2046204458cc18e8216d58d2ef983451501834605018347250183443501a205d58dc207e204c58fdd8d83465501834745018344650103447501a206dd8ec2046204458cc18e8216d58d2ef583459500834685008347a5008344b500a205d58dc207e2048346d5000344c500c58fdd8da206c18e8344e5000344f50093176300e297c2046204458cc18e8216d58d2ef183451500834605008344250003443500a205d58dc2046204458cc18d83465500834445000344650003457500a206c58e42046205418d558d02154d8d2aed03c5970183c5870183c6a70183c4b70122054d8dc206e204c58e558d83c5d70183c6c70183c4e70103c4f701a205d58dc2046204458cc18d82154d8d2afa03c5170183c5070183c6270183c4370122054d8dc206e204c58e558d83c5570183c6470183c4670103c47701a205d58dc2046204458cc18d82154d8d2af603c5970083c5870083c6a70083c4b70022054d8dc206e204c58e558d83c5d70083c6c70083c4e70003c4f700a205d58dc2046204458cc18d82154d8d2af203c5170083c5070083c6270083c4370022054d8dc206e204c58e558d83c5570083c6470083c4670083c77700a205d58dc204e207c58fdd8d82154d8d2aee01559307710b9304711315c103c4070083c60400fd14fd170505e308d4fe6363d40032833335d400aa939a8811a0b28813156700629503469501834685018347a5018344b5012206558ec207e204c58f5d8e8346d5018347c5018344e5010344f501a206dd8ec2046204458cc18e8216558e32f9034615018346050183472501834435012206558ec207e204c58f5d8e83465501834745018344650103447501a206dd8ec2046204458cc18e8216558e32f503469500834685008347a5008344b5002206558ec207e2048346d5000344c500c58fd18fa206c18e8344e5000344f50013166b006296c2046204458cc18e8216dd8e36f183461500834705008344250003443500a206dd8ec2046204458cc18e83475500834445000344650003457500a207c58f42046205418d5d8d0215558d2aed03459601834686018347a6018344b6012205558dc207e204c58f5d8d8346d6018347c6018344e6010344f601a206dd8ec2046204458cc18e8216558d2afa034516018346060183472601834436012205558dc207e204c58f5d8d83465601834746018344660103447601a206dd8ec2046204458cc18e8216558d2af603459600834686008347a6008344b6002205558dc207e204c58f5d8d8346d6008347c6008344e6000344f600a206dd8ec2046204458cc18e8216558d2af2034516008346060083472600834436002205558dc207e204c58f5d8d83465600834746008344660003467600a206dd8ec2046206458e558e0216518d2aee01551306710b9306711315c18347060083c40600fd167d160505e38897fe33b59700aa9363f597005a863a8b11a03a8613956800629583469501034785018347a5018344b501a206d98ec207e204c58fdd8e0347d5018347c5018344e5010344f50122075d8fc2046204458c418f0217d98e36f983461501034705018347250183443501a206d98ec207e204c58fdd8e0347550183474501834465010344750122075d8fc2046204458c418f0217d98e36f583469500034785008347a5008344b500a206d98ec207e2040347d5000344c500c58fd58f2207418f8344e5000344f50093166600e296c2046204458c418f02175d8f3af10347150083470500834425000344350022075d8fc2046204458c418f83475500834445000344650003457500a207c58f42046205418d5d8d0215598d2aed03c5960103c7860183c7a60183c4b6012205598dc207e204c58f5d8d03c7d60183c7c60183c4e60103c4f60122075d8fc2046204458c418f0217598d2afa03c5160103c7060183c7260183c436012205598dc207e204c58f5d8d03c7560183c7460183c4660103c4760122075d8fc2046204458c418f0217598d2af603c5960003c7860083c7a60083c4b6002205598dc207e204c58f5d8d03c7d60083c7c60083c4e60003c4f60022075d8fc2046204458c418f0217598d2af203c5160003c7060083c7260083c436002205598dc207e204c58f5d8d03c7560083c7460083c4660083c6760022075d8fc204e206c58ed98e8216558d2aee01559306710b130771130dc183c70600834407007d17fd160505e38897fe63e39700b28833b59700aa93468613156600629583469501034785018347a5018344b501a206d98ec207e204c58fdd8e0347d5018347c5018344e5010344f50122075d8fc2046204458c418f0217d98e36f983461501034705018347250183443501a206d98ec207e204c58fdd8e0347550183474501834465010344750122075d8fc2046204458c418f0217d98e36f583469500034785008347a5008344b500a206d98ec207e2040347d5000344c500c58fd58f2207418f8344e5000344f50093166b00e296c2046204458c418f02175d8f3af10347150083470500834425000344350022075d8fc2046204458c418f83475500834445000344650003457500a207c58f42046205418d5d8d0215598d2aed03c5960103c7860183c7a60183c4b6012205598dc207e204c58f5d8d03c7d60183c7c60183c4e60103c4f60122075d8fc2046204458c418f0217598d2afa03c5160103c7060183c7260183c436012205598dc207e204c58f5d8d03c7560183c7460183c4660103c4760122075d8fc2046204458c418f0217598d2af603c5960003c7860083c7a60083c4b6002205598dc207e204c58f5d8d03c7d60083c7c60083c4e60003c4f60022075d8fc2046204458c418f0217598d2af203c5160003c7060083c7260083c436002205598dc207e204c58f5d8d03c7560083c7460083c4660083c6760022075d8fc204e206c58ed98e8216558d2aee01559306710b130771130dc183c70600834407007d17fd160505e38897fe63f797002d4563f4a356850311a0328b13b513003375a8006319055a13146b00638f095ae3765b63b3048c0003c5990183c5890103c6a90183c6b90122054d8d4206e206558e518d83c5d90103c6c90183c6e90103c7f901a205d18dc2066207d98ed58d82154d8d2af903c5190183c5090103c6290183c6390122054d8d4206e206558e518d83c5590103c6490183c6690103c77901a205d18dc2066207d98ed58d82154d8d2af503c5990083c5890003c6a90083c6b90022054d8d4206e206558e518d83c5d90003c6c90083c6e90003c7f900a205d18dc2066207d98ed58d82154d8d2af103c5190083c5090003c6290083c6390022054d8d4206e206558e518d83c5590003c6490083c6690003c77900a205d18dc2066207d98ed58d82154d8d2aed03c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8d2afa03c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8d2af603c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8d2af203c5140083c5040003c6240083c6340022054d8d4206e206558e518d83c5540003c6440083c6640003c77400a205d18dc2066207d98ed58d82154d8d2aee01559305710b1306711301cd83c60500034706007d16fd150505e388e6fe63e5e63a4e89280a13060004e28597a00000e7804042130600046285a68597b00000e78020862c0a13060004268597a00000e780404093090c04280913060004e28597a00000e780003f0144568b1305fbff6370a414130871139308711b93156400ce954a76aa760a77ea6732fb36f73af33eef03c6950183c6850103c7a50183c7b5012206558e4207e2075d8f598e83c6d50103c7c50183c7e50183c4f501a206d98ec207e204c58fdd8e8216558e32fa03c6150183c6050103c7250183c735012206558e4207e2075d8f598e83c6550103c7450183c7650183c47501a206d98ec207e204c58fdd8e8216558e32f603c6950083c6850003c7a50083c7b5002206558e4207e2075d8f598e83c6d50003c7c50083c7e50083c4f500a206d98ec207e204c58fdd8e8216558e32f203c6150083c6050003c7250083c735002206558e4207e2075d8f598e83c6550003c7450083c7650083c57500a206d98ec207e205dd8dd58d8215d18d2eee81554686c28681cd0347060083c70600fd167d168505e308f7fe6366f7000504e319a4ec2a84637aa4162a8b93146500e2944a75aa750a76ea662afb2ef732f336ef03c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8d2afa03c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8d2af603c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8d2af203c5140083c5040003c6240083c6340022054d8d4206e20683c55400558e498e03c54400a20583c6640003c77400c98d1305fbffc2066207d98ed58d8215d18d2eee81551306711b9306711381cd0347060083c70600fd167d168505e308f7fee365f7ec131a64004e9a280a13060004d28597a00000e7808015130600045285a68597a00000e78060592c0a13060004268597a00000e78080130504a9b3930414002c0913060004628597a00000e7800012e3eb9a10b38a9a409a04269cca8963e47a016fe06f866fe0af80014593d81a0013966a00b304cc00e286130700fcb6873386e4000304060083850700238087002300b6000507850765f70505938404fc93860604e31b15fd134bfbff569b054585b46285d68597200000e780a0c40148fd3c6fe0cf816285d68597200000e78060d8e30305a46fd0fffa627c427a11a0568a13097113130d710be3784b076294280a13060004e28597a00000e7800007130600046285a28597a00000e780e04a2c0a13060004228597a00000e7800005930b0c04930afaffa80813060004e28597a00000e78080030144131564005e9583459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18d2ef983451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2ef583459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2ef183451500034605008346250003473500a205d18dc2066207d98ed58d034655008346450003476500034575002206558e42076205598d518d02154d8d2aed4675a6750676e6662afa2ef632f236ee01559305710b1306711305c183c60500034706007d16fd150505e388e6fe63f6e6000504e31754ed5684d685ae84637bb41213956400629583459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18d2ef983451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2ef583459500034685008346a5000347b500a205d18dc20662070346d500d98ecd8e8345c50022060347e5008347f5004d8e9385f4ff4207e2075d8f598e0216558e32f1034615008346050003472500834735002206558e4207e2075d8f598e83465500034745008347650003457500a206d98ec20762055d8d558d0215518d2aed46752676867666672afa32f636f23aee01556a86ca86e30105ee0347060083c70600fd167d160505e307f7fee376f7ec63ef845a62fc4ef066e852f863e79a5a814a8149014b814d26e43385844022f493156400de951a05338ca50093030008130300082eecae8b130871079302101033057c41135e650063775e0233b56d01b3b55901c98d3305b040137505f872952a8663e46d011e862a83b28389e513531500b303654063856d01639e5929a1aa630503148145130b81095e859308711b03469501834685010347a5018347b5012206558e4207e2075d8f598e8346d5010347c5018347e5010344f501a206d98ec2076204c18fdd8e8216558e32fb034615018346050103472501834735012206558e4207e2075d8f598e83465501034745018347650103447501a206d98ec2076204c18fdd8e8216558e32f703469500834685000347a5008347b5002206558e4207e2075d8f598e8346d5000347c5008347e5000344f500a206d98ec2076204c18fdd8e8216558e32f3034615008346050003472500834735002206558e4207e20783465500034445005d8f598ea206c18e03476500834775002300bb0085054207e2075d8fd98e8216558e32ef0156c686428715c283c7060003440700b3b48700a18f3334f000b3079040c18f7d17fd160506e5d311a0814713b6f7ff329b13050504e39665ec19a0130b8109930d810963925915638c03120145930a8111e2859308711b2380aa00050503c695fd83c685fd03c7a5fd83c7b5fd2206558e4207e2075d8f598e83c6d5fd03c7c5fd83c7e5fd83c4f5fda206d98ec207e204c58fdd8e8216558e32fb03c615fd83c605fd03c725fd83c735fd2206558e4207e2075d8f598e83c655fd03c745fd83c765fd83c475fda206d98ec207e204c58fdd8e8216558e32f703c695fc83c685fc03c7a5fc83c7b5fc2206558e4207e2075d8f598e83c6d5fc03c7c5fc83c7e5fc83c4f5fca206d98ec207e204c58fdd8e8216558e32f303c615fc83c605fc03c725fc83c735fc2206558e4207e2075d8f598e83c645fc03c755fc83c765fc83c475fc938505fc2207d98ec207e204c58fdd8e8216558e32ef0156c686428701ce83c70600034407007d17fd160506e38887fe33b68700b29ae31f75ec19a0930a8111930981113309bb4133853a416363a9002a896309090cf2e09ee49ae803c50d001a05b385ab00280b1306000497a00000e780e0a703ca090003c50d00934cfaff93956c00e2951a05de845e951306000497a00000e780a0a505456315a900ce8b6e8d99a87d1903c51d00138d1d001a053384a4001345faff136505f01a05629513060004a28597a00000e78040a203ca1900938b1900934cfaff93956c00e29513060004228597a00000e78040a07d19ea8dde89e31909fa13956c0062952c0b1306000497a00000e780609e930d1d0093891b001308710793021010a68b4663a663066e33c56d013335a0007d15337565001a05aa9b33c559013335a000b30570407d156d8d1a052a9ce3725ec263f86d0562840345fbff1309fbff1a05b384ab00130404fc280b13060004a68597a00000e780c097130600042685a28597a00000e780a0db2c0b13060004228597a00000e780c0954a8be3ee2dfb91a85e8463f8590503c5faff1389faff1345f5ff1a05b304ac00280b13060004a28597a00000e780c092130600042285a68597a00000e780a0d62c0b13060004268597a00000e780c09013040404ca8ae3ec29fb62653305a4401981a27aaa9aac08130600046274228597a00000e780408ec27463f99a0c139c6a00229c280a13060004a28597a00000e780808c130600042285e28597a00000e78060d02c0a13060004628597a00000e780808a33845441568963e38a0022897d1493090c04d54bc26c930d711363fe8a006275d6850276e68697d0ffffe780a07462f0a28a4e8c11a84e85a2856286e68697d0ffffe7802073627c2275a2653335b50013451500aae813d534003335a900134d150056f862fc827963e47a016fd02ff96fd08ff36285d68597100000e780809d6fd0cff35a85d68597a0ffffe780207e00005a85d285cdbf5685a685f5b72685ddb72285ddbf5d7186e4a2e026fc8505a5c12a8408659314150063e39500ae84914563e39500914497b5000083b5a5e8b3b5b400930640063386d402860509c918603305d5023af0894636f42af811a002f42800141097b0ffffe780e0a5a265426581cdfd55fe158505630ab50009ed9750ffffe780402c000008e004e4a6600664e2746161828062659750ffffe780002a0000130101dc233c1122233881222334912223302123233c312123384121368483c60600ba84b2892e8a2a89e5ce83c5040085e11385140097f5feff9385a5df1306000297a00000e78020b50125630905140a8597200000e78060ad0545230ca1100a852c0a05469760ffffe780e0aa230c41110a852c0a05469760ffffe780c0a90a8513060002ce859760ffffe780c0a8280aa28597000000e78080130a852c0a130600029760ffffe78000a7280aa68597000000e780c0110a852c0a130600029760ffffe78040a5280a8a851306800f97900000e780c0691304190002ea02e602e282fd280aac199770ffffe780605fac1913060002228597900000e7804067230009008330812303340123833481220339012283398121033a01211301012482801305140097f5feff9385a5d01306000297a00000e78020a683c5040001253366b50029e61385140097f5feff938565ce1306000297a00000e780e0a301250de9130610024a8581458330812303340123833481220339012283398121033a0121130101241793000067008351e31105ea05474a85d2854e86a68631a04a85d2854e86a28601478330812303340123833481220339012283398121033a012113010124170300006700e30f130101dc233c1122233881222334912223302123233c3121ae8483c505002a89d5c51384240093892402280097200000e780009309452300a11228000c1205469760ffffe7808090280013060002a2859760ffffe780808f280013060002ce859760ffffe780808e038514002300a11228000c1205469760ffffe780208d08122c001306800f97900000e780a05102ee02ea02e602e208120c029770ffffe78080470c02130600024a8597900000e780604f833081230334012383348122033901228339812113010124828093851400130600024a85833081230334012383348122033901228339812113010124179300006700234b130101da233c1124233881242334912423302125233c312323384123b68483c606002e892a84638a061403c5b40383c5a40303c6c40383c6d40322054d8d4206e206558e518d83c5f40303c6e40383c6040483c71404a205d18dc206e207dd8ed58d82154d8daaea03c5340383c5240303c6440383c6540322054d8d4206e206558e518d83c5740303c6640383c6840383c79403a205d18dc206e207dd8ed58d82154d8daae603c5b40283c5a40203c6c40283c6d40222054d8d4206e206558e518d83c5f40203c6e40283c6040383c71403a205d18dc206e207dd8ed58d82154d8daae203c5340283c5240203c6440283c6540222054d8d4206e20683c57402558e518d03c66402a20583c6840283c794024d8e93852400c206e207dd8e558e0216518d2afe05c3131589036d91301a329503060500937679000547b316d700558e2300c500130524001306000297900000e780c035130524022c1a1306000297900000e780a034038514000525a300a40005452300a4007da8b289850402ec02e802e402e005c3131589036d918a852e95830505001376790085463396c600d18d2300b500130a2400081097100000e780a06b230c211308102c1a054605499750ffffe7802069081013060002ce859750ffffe7802068081013060002a6859750ffffe7802067281a0c101306800f97900000e780a02b02fa02f602f202ee281a2c0a9770ffffe78080212c0a13060002528597900000e7806029130524028a851306000297900000e7804028a3002401230024018330812503340125833481240339012483398123033a0123130101268280157186eda2e9a6e5cae14efd52f956f55af15eed62e966e5328a7d16637ab63c2e89637aba3aaa89930a7102130b7108930b7108130c71065284050a93146400ce9403c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8d2ae103c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8daafc03c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8daaf803c5140083c5040003c6240083c6340022054d8d4206e206558e518d83c5540003c6440083c6640003c77400a205d18dc2066207d98ed58d82154d8daaf403c594fd83c584fd03c6a4fd83c6b4fd22054d8d4206e206558e518d83c5d4fd03c6c4fd83c6e4fd03c7f4fda205d18dc2066207d98ed58d82154d8d2af003c514fd83c504fd03c624fd83c634fd22054d8d4206e206558e518d83c554fd03c644fd83c664fd03c774fda205d18dc2066207d98ed58d82154d8d2aec03c594fc83c584fc03c6a4fc83c6b4fc22054d8d4206e206558e518d83c5d4fc03c6c4fc83c6e4fc03c7f4fca205d18dc2066207d98ed58d82154d8d2ae803c514fc83c504fc03c624fc83c634fc22054d8d4206e20683c554fc558e518d03c644fca20583c664fc03c774fcd18d938c04fcc2066207d98ed58d82154d8d2ae40155da855686630b051883c60500034706007d16fd150505e387e6fe63f0e618280013060004a68597900000e78080ff130600042685e68597900000e78080fe7d14630504147d1493146400ce940275e2654266a266aaf0aeecb2e8b6e403c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8d2ae103c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8daafc03c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8daaf803c5140083c5040003c6240083c6340022054d8d4206e206558e518d83c5540003c6440083c6640003c77400a205d18dc2066207d98ed58d82154d8daaf40155e2855e8605c983c60500034706007d16fd150505e388e6fe63fee600130600046685a68597900000e78040eaa68ce31004ecce8c2c0013060004668597900000e780c0e8e3132ac7ee604e64ae640e69ea794a7aaa7a0a7bea6b4a6caa6c2d61828017e5feff130585599305e0029790ffffe78000580000317106fd22f926f54af14eed52e956e55ae1defce2f8e6f4eaf02e89aa8993da1500130bf103930bf101130cf103930cf101fd1a13961a00130816006377284956850906637f262193166800ce9603c7960183c7860183c4a60103c4b60122075d8fc2046204458c418f83c7d60183c4c60103c4e60183c5f601a207c58f4204e205c18ddd8d8215d98d2eec83c5160103c7060183c7260183c43601a205d98dc207e204c58fdd8d03c7560183c7460183c4660103c4760122075d8fc2046204458c418f0217d98d2ee883c5960003c7860083c7a60083c4b600a205d98dc207e20403c7d60003c4c600c58fdd8d2207418f83c7e60083c4f6001a064e96c207e204c58f5d8f0217d98d2ee483c5160003c7060083c7260083c43600a205d98dc207e204c58fdd8d03c7560083c7460083c4660083c6760022075d8fc204e206c58ed98e8216d58d2ee083459601834686010347a6018347b601a205d58d4207e2075d8fd98d8346d6010347c6018347e6018344f601a206d98ec207e204c58fdd8e8216d58d2efc83451601834606010347260183473601a205d58d4207e2075d8fd98d83465601034746018347660183447601a206d98ec207e204c58fdd8e8216d58d2ef883459600834686000347a6008347b600a205d58d4207e2075d8fd98d8346d6000347c6008347e6008344f600a206d98ec207e204c58fdd8e8216d58d2ef483451600834606000347260083473600a205d58d4207e2075d8fd98d83465600034746008347660003467600a206d98ec20762065d8e558e0216d18d2ef00156de865a8719ce83c70600834407007d17fd160506e38897fe33ba970021a0428a19a0014a429a6379257763742a771a053384a90093146a00ce9403459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8d2aec0345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8d2ae803459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8d2ae40345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8d2ae003c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8d2afc03c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8d2af803c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8d2af403c5140083c5040003c6240083c6340022054d8d4206e206558e518d83c5540003c6440083c6640003c77400a205d18dc2066207d98ed58d82154d8d2af00155e685628639c983c60500034706007d16fd150505e388e6fe63f1e604081013060004a28597900000e780c09b130600042285a68597900000e780a0df0c1013060004268597900000e780c09913161a00130816005285e36e28b7e3940ab6130bf103930bf101130cf103930cf101094dca8afd1a63fb2a4f13946a004e94081013060004ce8597900000e780a095130600044e85a28597900000e78080d90c1013060004228597900000e780a09363ebaa490146014505480906637f562193166800ce9603c7960183c7860183c4a60103c4b60122075d8fc2046204458c418f83c7d60183c4c60103c4e60183c5f601a207c58f4204e205c18ddd8d8215d98d2eec83c5160103c7060183c7260183c43601a205d98dc207e204c58fdd8d03c7560183c7460183c4660103c4760122075d8fc2046204458c418f0217d98d2ee883c5960003c7860083c7a60083c4b600a205d98dc207e20403c7d60003c4c600c58fdd8d2207418f83c7e60083c4f6001a064e96c207e204c58f5d8f0217d98d2ee483c5160003c7060083c7260083c43600a205d98dc207e204c58fdd8d03c7560083c7460083c4660083c6760022075d8fc204e206c58ed98e8216d58d2ee083459601834686010347a6018347b601a205d58d4207e2075d8fd98d8346d6010347c6018347e6018344f601a206d98ec207e204c58fdd8e8216d58d2efc83451601834606010347260183473601a205d58d4207e2075d8fd98d83465601034746018347660183447601a206d98ec207e204c58fdd8e8216d58d2ef883459600834686000347a6008347b600a205d58d4207e2075d8fd98d8346d6000347c6008347e6008344f600a206d98ec207e204c58fdd8e8216d58d2ef483451600834606000347260083473600a205d58d4207e2075d8fd98d83465600034746008347660003467600a206d98ec20762065d8e558e0216d18d2ef00156de865a8719ce83c70600834407007d17fd160506e38897fe33ba970021a0428a19a0014a429a63715529637e5a271a053384a90093146a00ce9403459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8d2aec0345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8d2ae803459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8d2ae40345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8d2ae003c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8d2afc03c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8d2af803c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8d2af403c5140083c5040003c6240083c6340022054d8d4206e206558e518d83c5540003c6440083c6640003c77400a205d18dc2066207d98ed58d82154d8d2af00155e6856286e30405b883c60500034706007d16fd150505e387e6fee3f9e6b6081013060004a28597800000e780404d130600042285a68597900000e78020910c1013060004268597800000e780404b13161a00130816005285e36d58b705beea704a74aa740a79ea694a6aaa6a0a6be67b467ca67c067d296182805285d68529a0528511a05685ca859790ffffe780c0430000757106e522e1a6fccaf8cef4d2f0d6ecdae8dee4ae89fd1513d61500d18d13d62500d18d13d64500d18d13d68500d18d13d60501d18d13d60502d18d93c5f5ff17a60000033626ae97a6000083b626ae13d71500798e918d33f6d5008981f58db29517a60000033606ad97a6000083b606ad13d74500ba95f18db385d502e1917d56b35ab600850a638a0a0a2a8913d519007999fd1a130bf5ff13d529001e054a95130405fc8d44ce8b63723b091395db0033457501935575002d8d93151501b3cba50033f55b01b3353501fd15b3f535010d8d637e35051a05330aa900280013060004a28597800000e7802038130600042285d28597800000e780007c2c0013060004528597800000e7802036050bfd1413040404d1f8aa600a64e6744679a679067ae66a466ba66b496182805a85ce859790ffffe7800030000017e5feff1305e5a3f1459790ffffe78080a40000557186e5a2e126fd4af94ef552f156ed5ae95ee562e1e6fceaf8eef42e8c2a89014b930b7104930c710213bd2503954d854463f384238545139564004a9503469501834685010347a5018347b5012206558e4207e2075d8f598e8346d5010347c5018347e5010344f501a206d98ec2076204c18fdd8e8216558e32f0034615018346050103472501834735012206558e4207e2075d8f598e83465501034745018347650103447501a206d98ec2076204c18fdd8e8216558e32ec03469500834685000347a5008347b5002206558e4207e2075d8f598e8346d5000347c5008347e5000344f500a206d98ec2076204c18fdd8e8216558e32e8034615008346050003472500834735002206558e4207e2075d8f598e83465500034745008347650003447500a206d98ec2076204c18fdd8e8216558e32e4034695fd834685fd0347a5fd8347b5fd2206558e4207e2075d8f598e8346d5fd0347c5fd8347e5fd0344f5fda206d98ec2076204c18fdd8e8216558eb2e0034615fd834605fd034725fd834735fd2206558e4207e2075d8f598e834655fd034745fd834765fd034475fda206d98ec2076204c18fdd8e8216558e32fc034695fc834685fc0347a5fc8347b5fc2206558e4207e2075d8f598e8346d5fc0347c5fc8347e5fc0344f5fca206d98ec2076204c18fdd8e8216558e32f8034615fc834605fc034725fc834735fc2206558e4207e2075d8f598e834655fc034745fc834765fc034575fca206d98ec20762055d8d558d0215518d2af401556686de8601cd0347060083c70600fd167d160505e308f7fe6369f7008504b3b58401e39384df51a0814533c58401133515003366ad003dea9389f4ff63f789098589d1c5139a69004a9a939a6400ca9a281013060004d28597800000e7800009130600045285d68597800000e78000082c1013060004568597800000e78000070545637f95004a85a6854e8697f0ffffe78060e04a85a68597000000e7804004050be310bbd7014511a00545ae600e64ea744a79aa790a7aea6a4a6baa6b0a6ce67c467da67d696182804e8511a02685e2859790ffffe78000fe0000317106fd22f926f54af14eed52e956e55ae12e89aa840345950583c5840503c6a40583c6b40522054d8d4206e206558e518d83c5d40503c6c40583c6e40503c7f405a205d18dc2066207d98ed58d82154d8daafc03c5140583c5040503c6240583c6340522054d8d4206e206558e518d83c5540503c6440583c6640503c77405a205d18dc2066207d98ed58d82154d8daaf803c5940483c5840403c6a40483c6b40422054d8d4206e206558e518d83c5d40403c6c40483c6e40403c7f404a205d18dc2066207d98ed58d82154d8daaf403c5140483c5040403c6240483c6340422054d8d4206e206558e518d83c5540403c6440483c6640403c77404a205d18dc2066207d98ed58d82154d8daaf003c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8d2aec03c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8d2ae803c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8d2ae403c5140083c5040003c6240083c6340022054d8d4206e20683c55400558e518d03c64400a20583c6640003c77400d18d93890404c2066207d98ed58d82154d8d2ae01305f10181551306f1076380051a83460600034705007d157d168505e387e6fe63f5e6180a8513060004a68597800000e78060dd130600042685ce8597800000e78060dc0d45636aa914130af107894a130bf10513946a00269403459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8daaec0345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8daae803459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8daae40345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8daae06265c26522668266aafcaef8b2f4b6f00155da8552860dc983c60500034706007d16fd150505e388e6fe63ffe600850a130504fc13060004a28597800000e78060c7a289e39f2aeb8a85130600044e8597800000e78000c6ea704a74aa740a79ea694a6aaa6a0a6b29618280257106ef22eb26e74ae32a8484004800130901031306c002814597800000e780c0b5130680132685814597800000e780c0b417d5feff9305550741464a8597800000e78060c0370501011b0505022ac082fe8a8522859740ffffe78000e4fa605a64ba641a691d6182805d7186e4a2e026fc8505a5c12a8408659314150063e39500ae84914563e3950091449795000083b52529b3b5b400930600053386d4028e0509c918603305d5023af0a14636f42af811a002f4280014109790ffffe780e0e3a265426581cdfd55fe158505630ab50009ed9730ffffe780406a000008e004e4a6600664e2746161828062659730ffffe780006800005d7186e4a2e026fc4af8ae84806590612a892800a2859770ffffe78080400345810001c9426505c59780ffffe7806041000005040dc49305910080e4130519001306000297800000e78080b005452300a900a6600664e27442796161828017d5feff13050520f1459780ffffe780a02000000e0597d5feff938525962e950c6105458285094582800d458280114582809780ffffe780e03a0000106195456316b60003058500050582800c65328517030000670043fc130101d32334112c2330812c233c912a2338212b2334312b2330412bb2842e842a8902f002ec02e802e4930901164812130a01151306c002814597800000e780e098130680134e85814597800000e780e09717d5feff930575ea4146528597800000e78080a3370501011b0505022320a112233c012828100c129740ffffe780e0c62810a28526869740ffffe78060db08122c101306800f97800000e780e09f08122c009760ffffe78040962c00130600024a8597800000e780209e8330812c0334012c8334812b0339012b8339812a033a012a1301012d8280317106fd22f926f54af14eed52e993070002631cf61eba89368a2a8903c5950103c6850183c6a50103c7b5012205518dc2066207d98e558d03c6d50183c6c50103c7e50183c7f5012206558e4207e2075d8f598e0216518d2aec03c5150103c6050183c6250103c735012205518dc2066207d98e558d03c6550183c6450103c7650183c775012206558e4207e2075d8f598e0216518d2ae803c5950003c6850083c6a50003c7b5002205518dc2066207d98e558d03c6d50083c6c50003c7e50083c7f5002206558e4207e2075d8f598e0216518d2ae403c5150003c6050083c6250003c735002205518dc2066207d98e558d03c6550083c6450003c7650083c575002206558e4207e205d98dd18d82154d8d2ae088009770ffffe78040c6a8188a859770ffffe78000b3266511c506659730ffffe780e0392a658a6566762afc2ef832f40305710783056107e664034651072303a102a20503452107d18d2312b10283451107220503463107830641074d8d06744206e206558e518d2ad0a818d2854e869770ffffe780e0b111c426859730ffffe780e0332275e6754276aae062758a66b2e42a66aae8aeecb6f0b2f405452308a106130511070c101d4697700000e780e07fa8188c009770ffffe78020c3880097000000e780600566742a664a85a28597000000e78020d40a6511c522859730ffffe780c02dea704a74aa740a79ea694a6a2961828017d5feff130525f197d5feff9386c5f39305b00290009780ffffe78020070000411106e422e02a84086511c508609730ffffe7806029087009c9086ca260026441011733ffff67002328a260026441018280697106f622f226ee4aea4ee652e2d6fddaf9def5e2f1e6ed2e8a2a89014481490d45aae082e49304110501163335c00093b51500b36ab500130b1108894b7d5c88088c009790ffffe780a051034501056309751f6301051003c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8d2ae903c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8d2ae503c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8d2ae103c5140083c5040003c6240083c6340022054d8d4206e206558e518d83c5540003c6440083c6640003c77400a205d18dc2066207d98ed58d82154d8daafc63890a00dda002e902e502e182fc639e0a0ca81813060002d28597800000e780e0a1012579e1639a091628110d46a2859770ffffe780e0fa2a7559c96a75ca752a76aae9aee5b2e1a8188c019790ffffe78020220305eb008305db000346cb00e6792303a10aa205d18d2312b10a03459b0083458b000346ab008306bb0022054d8d4206e206558e518d2ad103451b0083450b0003462b0083463b0022054d8d4206e20683455b00558e518d03464b00a20583466b0003477b00d18d834c0108c2066207d98ed58d82154d8d2aed11a081496a658a550316410a8306610a2af82edc231ec102230fd102630e8409050401b5638609060305e1038315c1036256c2762307a1022316b10232d436f0130511010c103d4697700000e780a04f4ee423089101a8182c0005469790ffffe78080d6667535c92a658a656676aaf0aeecb2e888089790ffffe78080f12334a9004e859790ffffe78060a4014531a01305a005a300a90005452300a900b2701274f2645269b269126aee7a4e7bae7b0e7cee6c5561828017d5feff1305c5b9f1459780ffffe78060ba000017d5feff130585ec9305b002edb717d5feff130585bc97c5feff9386253c9305b00290089780ffffe78080d20000497186f6a2f2a6eecaeacee6d2e256fe5afa5ef662f266ee6aea6ee62e842ae0814a014d0149014b0945aaf882fc93041108bd497d5a2ee408018c1897000000e780008c03450108630b052803c5940183c5840103c6a40183c6b40122054d8d4206e206558e518d83c5d40103c6c40183c6e40103c7f401a205d18dc2066207d98ed58d82154d8daae103c5140183c5040103c6240183c6340122054d8d4206e206558e518d83c5540103c6440183c6640103c77401a205d18dc2066207d98ed58d82154d8d2afd03c5940083c5840003c6a40083c6b40022054d8d4206e206558e518d83c5d40003c6c40083c6e40003c7f400a205d18dc2066207d98ed58d82154d8d2af903c5140083c5040003c6240083c6340022054d8d4206e206558e518d83c5540003c6440083c6640003c77400a205d18dc2066207d98ed58d82154d8d2af5281113060002a28597700000e780407201256310051888190946d6859770ffffe78060cbce7b638a0b1e126c6e7563fc8915aae8eaec414581459780ffffe78060642a842e8b4146de8597700000e780a02b83458400834994000349a400834db4000346c400034dd4008347e400034af400834c04000347140083432400834634000348440003435400834864008342740063050b04228542f0468416fc6aec1a8d4ae81e896ef4b68dcee0ba89b2e452f83e8a2e8b9730ffffe78000d6da85d287427a26664e878669ee86a27dca8342696a83626de272a28802786665631e0514a20933e5b9004209e20db3e52d014d8d220db365cd0013960701620a3366ca00d18d8215b3eda50013158700336595019395030113968601d18d4d8d93158300b3e505011396080193968201558ed18d8215b3eca50013040cff93890b01228581459780ffffe780c0532a8c2e8bce85228697700000e780001be2f9dafd22e2a8098c199790ffffe780c0df8c1188618c65014b6e6daaf0aef405492264bd497d5a466511c55e859730ffffe780c0c8638a4a07850ab1bb3365690119cd630d0d0226758675026608f20cee233096012334b6012338a6013da01305500382652380a50023b80500630f0d006a859780ffffe780c06b01a81305200382652380a50023b80500b6701674f6645669b669166af27a527bb27b127cf26c526db26d7561828017d5feff13050581f1459780ffffe780a081000017d5feff1305a58497d5feff938645899305b002b0099780ffffe780a09a000017d5feff130575b493059002e9b7097186fea2faa6f6caf2ceeed2ead6e6dae25efe62fa66f66af26eeeb289ae842ae4014b014d0149814b32e102e5130411093d4afd5a32ec2ee808090c0197f0ffffe780205303450109630c052803459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8daae90345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8daae503459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8daae10345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8d2afd281913060002a68597700000e78060390125631105180802da854e869770ffffe7808092126c630b0c1ed26c3265637d9a15aaf0eaf4414581459780ffffe780802baa84ae8b4146e28597700000e780c0f283c5840003ca940003c9a40083c9b40003c6c40083cdd40083c7e40083caf40003cd040003c7140083c3240083c6340003c8440003c3540083c8640083c2740063850b042685c28bc684d6e016f86ef49a8d4af01e89b6e4d2e83a8ab2ec4efcbe89ae8a9730ffffe780209dd685ce87e27966665287466aa666ca8302796e83a27dc272866aa6885e882675631f0514220a3365ba004209e209b3e529014d8da20db3e5cd0013960701e20a33e6ca00d18d82154d8daaf4131587003365a5019395030113968601d18d4d8d93158300b3e505011396080193968201558ed18d8215b3eda50093840cff130a0c01268581459780ffffe780e01aaa8cae8bd285268697700000e78020e266e25ee626eaa8110c029790ffffe780e0a68c1988618c65814b2e7daaf8aefc0549e269c2643d4afd5a067511c562859730ffffe780c08f630a5b07050ba9bb3365790119cd630d0d026675c675226608f20cee2330b601267508e62338a6013da013055003a2652380a50023b80500630f0d006a859780ffffe780c03201a813052003a2652380a50023b80500f6705674b6741679f669566ab66a166bf27b527cb27c127df26d1961828017c5feff13050548f1459770ffffe780a048000017c5feff1305a54b97c5feff938645509305b002b0119770ffffe780a061000017c5feff1305057e9305c002e9b7097186fea2faa6f6caf2ceeed2ead6e6dae25efe62fa66f66af26eeeae892ae4014b814a214a52e802ec02f005452af402f8130d9103930d110b0944fd5428182c109790ffffe78080ae034581036309853475cd03459d0183458d010346ad018346bd0122054d8d4206e206558e518d8345dd010346cd018346ed010347fd01a205d18dc2066207d98ed58d82154d8daae503451d0183450d0103462d0183463d0122054d8d4206e206558e518d83455d0103464d0183466d0103477d01a205d18dc2066207d98ed58d82154d8daae103459d0083458d000346ad008346bd0022054d8d4206e206558e518d8345dd000346cd008346ed000347fd00a205d18dc2066207d98ed58d82154d8d2afd03451d0083450d0003462d0083463d0022054d8d4206e206558e518d83455d0003464d0083466d0003477d00a205d18dc2066207d98ed58d82154d8d2af929a082e582e102fd02f9081913060002ce8597700000e78060ff01256318052208190546da859760ffffe780c0480345010b6311052603c59d0183c58d0103c6ad0183c6bd0122054d8d4206e206558e518d83c5dd0103c6cd0183c6ed0103c7fd01a205d18dc2066207d98ed58d82154d8daafc03c51d0183c50d0103c62d0183c63d0122054d8d4206e206558e518d83c55d0103c64d0183c66d0103c77d01a205d18dc2066207d98ed58d82154d8daaf803c59d0083c58d0003c6ad0083c6bd0022054d8d4206e206558e518d83c5dd0003c6cd0083c6ed0003c7fd00a205d18dc2066207d98ed58d82154d8daaf403c51d0083c50d0003c62d0083c63d0022054d8d4206e206558e518d83c55d0003c64d0083c66d0003c77d00a205d18dc2066207d98ed58d82154d8daaf008190546da859760ffffe780a047ca7b63870b168e653d456378b51a6a79138405ff138c0b01228581459780ffffe78040e0aa84ae8ce285228697700000e78080a726f966fda2e108010c199780ffffe780406c28090c019730ffffe780609608020c010d469780ffffe780e02c1265630305125265b2651266aae12efd32f908020c199780ffffe78000575265d145631cb510126451468809a28597700000e78060a13265fd5411c522859720ffffe78080510675a67546762af92efdb2e16675aa750a76ea666267aae5a8110ce910e514e1639aea000808d68597f0ffffe780c0df827a426a0944130500053385aa0252950c191306000597700000e780809b0a65850a56f09780ffffe78020f3630709005e859720ffffe780e04a630a9b02050b45b10275e2654266a26688ea8ce690e2f6705674b6741679f669566ab66a166bf27b527cb27c127df26d1961828017c5feff13052507f1459770ffffe780c007000017c5feff1305c50a97c5feff9386650f9305b002901089a017c5feff1305450997c5feff9386e50d9305b00210022da017c5feff1305c50797c5feff9386658709a817c5feff1305a50697c5feff938645099305b00210199770ffffe780a01c000041459780ffffe780208b0000757106e522e1a6fccaf8cef4d2f02a89814432e402e81304910181153335b00093351900b369b500094a28082c009780ffffe780e06a0345810165d9630c451303459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8daaec0345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8daae803459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8daae40345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8daae0e39909ee880013060002ca8597700000e78020bc0125e31e05ec93f4f40f850413f5f40fe30795ec17c5feff130505e9f1459770ffffe780a0e900002685aa600a64e6744679a679067a49618280517186f5a2f1a6edcae9cee5d2e156fd5af95ef562f166ed6ae96ee5b2892e8a2ae0014b814a32ec02f013049102894d7d5928102c089780ffffe7800052034581026300b51b75cd03459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8daaf40345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8daaf003459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8daaec0345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8daae829a082f482f082ec82e8880813060002d28597700000e780e0a2012519c1d684a5a88808da854e869760ffffe780e0fbc66b63820b0c666d8674268581459780ffffe7806095aa8c2e8cde85268697600000e780a05ce6e8e2eca6f088188c089780ffffe7806021ac1888618c65c674aae8aeec63870a0056859780ffffe78060b26665c6652ae82ee463070d005e859720ffffe780a00963052b05050ba68a89bd63890a004265a265026608ea32850ce639a01305b00682652384a5002e8523305501ae700e74ee644e69ae690e6aea7a4a7baa7b0a7cea6c4a6daa6d6d61828017c5feff130585c4f1459770ffffe78020c5000017c5feff130525c897c5feff9386c5cc9305b00290189770ffffe78020de00001d7186eca2e8a6e4cae02a84081097000000e780c0d98274a1c40309810293059102130511013d4697600000e780a04d26e42308210108102c000d469780ffffe78080d402750dc94275a275027608e80ce410e026859780ffffe78040a339a0030581022304a40023300400e6604664a66406692561828017c5feff1305a5be97b5feff9386453e9305b0021306f1039770ffffe78080d40000357106ed22e926e5aa85a8100d4697000000e78020d0267461c88304010793051107130511013d4697600000e780004422e423089100a8102c0011469780ffffe780e0ca26754dcd6675c67526762af82ef432f0a8100c1001469780ffffe78000c926755dc56675c6752676aae4aee032fc88082c1809469780ffffe78020c7466545c50675e6654666aafcaef8b2f4231201088808ac105001894689449780ffffe780809a0345010541ed6665631b950a8314410826759780ffffe780809362759780ffffe780e09202759780ffffe780409222859780ffffe780a091014501469b95040131a003450107814522050546d18d4d8dea604a64aa640d61828017c5feff130585ac97b5feff9386252c09a817c5feff130565ab97b5feff9386052b9305b00290080da817c5feff1305e5a997b5feff938685299305b002b01029a817c5feff130565a897c5feff938605809305b002130671089770ffffe78040be000017c5feff1305c591b9459770ffffe78000a20000517186f5a2f1a6edcae9cee5d2e156fd5af95ef562f166ed6ae96ee5b2892e8a2ae0014b814a32ec02f013049102894d7d5928102c089780ffffe780800b034581026300b51b75cd03459401834584010346a4018346b40122054d8d4206e206558e518d8345d4010346c4018346e4010347f401a205d18dc2066207d98ed58d82154d8daaf40345140183450401034624018346340122054d8d4206e206558e518d83455401034644018346640103477401a205d18dc2066207d98ed58d82154d8daaf003459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8daaec0345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8daae829a082f482f082ec82e8880813060002d28597600000e780605c012519c1d684a5a88808da854e869760ffffe78060b5c66b638a0b0a666d8674268581459770ffffe780e04eaa8c2e8cde85268697600000e7802016e6e8e2eca6f088188c089780ffffe780e0daac1888618c65c674aae8aeec63870a0056859770ffffe780e06b6665c6652ae82ee463070d005e859720ffffe78020c3630d2b03050ba68a89bd63820a064265a265026608ea0ce623305601ae700e74ee644e69ae690e6aea7a4a7baa7b0a7cea6c4a6daa6d6d61828017b5feff1305057ff1459760ffffe780a07f000017c5feff1305a58297c5feff938645879305b00290189770ffffe780a098000017b5feff1305e5789305b002e9b7130101ce233c1130233881302334913023302131233c312f2338412f2334512f2330612f233c712d2338812d2334912d2330a12d233cb12b3a8a3684328bae892a891305000285459720ffffe780e0b56306056eaa8413060002814597600000e78020f7514585459720ffffe780e0b36309056c2a8c5146814597600000e78040f51305000281459770ffffe7800039aa8bae8a13060002d28597600000e780200026859720ffffe780a0b00345140183450401034624018306340122054d8d4206e206558e518daac803459400834584000346a4008346b40022054d8d4206e206558e518d8345d4000346c4008346e4000347f400a205d18dc2066207d98ed58d82154d8daae40345140083450400034624008346340022054d8d4206e206558e518d83455400034644008346640003477400a205d18dc2066207d98ed58d82154d8daae0130a0105930c8104514581459770ffffe780602c2afeaee282e693041104281a8c0026869770ffffe780601113042104281aa68522869770ffffe780401093043104281aa28526869770ffffe780200fc000281aa68522869770ffffe780200e93045104281aa28526869770ffffe780000d13046104281aa68522869770ffffe780e00b93047104281aa28526869770ffffe780c00a281aa68566869770ffffe780e00913049104281ae68522869770ffffe780c0089304a104281aa28526869770ffffe780a0071304b104281aa68522869770ffffe7808006e400281aa28526869770ffffe78080051304d104281aa68522869770ffffe78060049304e104281aa28526869770ffffe78040031304f104281aa68522869770ffffe7802002281aa28552869770ffffe780400113041105281ad28522869770ffffe780200093042105281aa28526869770ffffe78000ff13043105281aa68522869770ffffe780e0fdd008281aa2859770ffffe78000fdf27c966d366a62859720ffffe780e08e1304ca02636e4445228581459770ffffe78040142afeaee282e64145a1459720ffffe780008c630c05442a8c31452330ac001305c0022334ac00a2c0d000281a8c009770ffffe78060f78944130d410462840860aac0281a8c006a869770ffffe780c0f5fd142104edf462859720ffffe780a08713860b02281ade859770ffffe780c0f333864c01281ae6859770ffffe780c0f2727a166d366c63870a005e859720ffffe780608463870d0066859720ffffe78080835a8581459770ffffe78060092a84ae8ace855a8697600000e780a0d013050002631aab3a03056400230fa112030554008345440022054d8d231ea1120345140083450400034624008306340022054d8d4206e206558e518d232ca1120345840083457400034694008346a40022054d8d4206e206558e518d8345c4000346b4008346d4000347e400a205d18dc2066207d98ed58d8215b3e9a500034504018345f400034614018346240122054d8d4206e206558e518d83454401034634018346540103476401a205d18dc2066207d98ed58d8215b3eba5000345840183457401034694018346a40122054d8d4206e206558e518d8345c4010346b4018346d4010347e401a205d18dc2066207d98e034bf401d58d8215b3e4a50063870a0022859710ffffe78000710305e1138315c113032681132303a1042312b104b2c0a303310513d589032307a10413d50903a306a10413d589022306a10413d50902a305a10413d589012305a10413d50901a304a10413d589002304a104a307710513d58b03230ba10413d50b03a30aa10413d58b02230aa10413d50b02a309a10413d58b012309a10413d50b01a308a10413d58b002308a104a30b910413d58403230fa10413d50403a30ea10413d58402230ea10413d50402a30da10413d58401230da10413d50401a30ca104a180230c9104a30f6105281a9750ffffe78060ee08108c009750ffffe78020db166511c572759710ffffe78000624275a27502762aec2ee832e40305f1168305e11656640346d1162303a100a2050345a116d18d2312b1008345911622050346b1168306c1164d8df6644206e206558e518d2ac00810d28562869750ffffe78000da91c422859710ffffe780005c2265827542662afe6265a276b2e24276aae6aeeab6eeb2f205452304a116130591168a851d4697600000e78000a828002c1a9750ffffe78040eb281a97e0ffffe780802d02fc02f802f402f0a01a681aa4121306c002814597600000e7800098130680132285814597600000e780009717b5feff930595e94146268597600000e780a0a2370501011b050502232ca1122338012a88002c1a9720ffffe78000c6226462668800a2859720ffffe78060da281a8c001306800f97600000e780e09e281a0c109740ffffe78040950c10130600024a8597600000e780209d426511c522859710ffffe780604d63070d0052859710ffffe780804c833081310334013183348130033901308339812f033a012f833a812e033b012e833b812d033c012d833c812c033d012c833d812b13010132828017b5feff1305658ff1459760ffffe780000900001305000221a0514511a041459710ffffe780e047000017b5feff1305a50a97b5feff938645119305b002301a9760ffffe780a0200000130101dd2334112223308122233c91202e84aa8402f002ec02e802e4281097e0ffffe78080cc22f228100c1221469720ffffe78040ca08122c101306800f97600000e780c08e08122c009740ffffe78020852c0013060002268597600000e780008d833081220334012283348121130101238280130101812334117e2330817e233c917c2338217d2334317d2330417d233c517b2338617b2334717b2330817b233c91792338a1792334b179357136ec32e42ee82a842338014623340146a80813068002814597500000e78060790335014683358146033601472ae12ee5086032e902f10c683336a00014643307c040f98d32f502f92afdb6e1b2e582e9aaedb6f1aef5130da122930ba124854d930a400828119770ffffe780606819e16f2090222a8493040501233c0178233801782334017823300178881697e0ffffe780c0ba88165146a6859720ffffe780a0b8130501468c161306800f97500000e780007d13050146930501789730ffffe7802073033581798335017903368178833601782ae62ee2b2fdb6f9033b0400033c84002af62ef232ee36ea233c0178233801782334017823300178881697e0ffffe780a0b3233481472330614788169305014641469720ffffe780e0b0130501468c161306800f97500000e780407513050146930501789730ffffe780606b930501781306000213041113228597500000e780e0722308011217b5feff930565de13060002228597600000e780c0b3012521c1327592757266d2664a6a2334a1282330b128233cc1262338d12663080a046a648c1c52859770ffffe7808077ae842dcd41c48e04d29403ba04227d14d5b74a64e30a04386a65b384ad400c0a22859770ffffe780e07463000518e38db4378e05a29503b405228504cdb7833981278334012803398128033401279770ffffe780e05b233805208545231db52000e12334350104e9233c250123348517233065172ae902ed6f00f0329204d29423b4841723b064176f001032033d812783350128833c81280359aa21833b01272d456379a91293891400139454005294939a44006375391d2300740113d58b03a303a40013d50b032303a40013d58b02a302a40013d50b022302a40013d58b01a301a40013d50b012301a40013d58b00a300a4002304a40113558d03a307a40013550d032307a40013558d02a306a40013550d022306a40013558d01a305a40013550d012305a40013558d00a304a4002308b40013d58503a30ba40013d50503230ba40013d58502a30aa40013d50502230aa40013d58501a309a40013d505012309a40013d58500a308a400230c940113d58c03a30fa40013d50c03230fa40013d58c02a30ea40013d50c02230ea40013d58c01a30da40013d50c01230da40013d58c00a30ca400f5aa2300015a639ab40323308136233401362338b136130501468c161306015a9770ffffe78040616f20206f854d1545aee463f2a41e1149e5aa8e05a29503b5052299c8b30590400356a5210e06329503350522fd15edf98355a521fd152338a164233c01642330b16613050146930501651306015a9770ffffe780e05b0335814783350147233ca17803368146833601462338b178033501492334c1782330d1780339014a8355a521833481492a846374b9006f20004e0334052119e06f20204d035985218355a42185042285e375b9fe6f20204c139559005295b304994013965400d6e8ae8aa28597600000e780808913d58b03a303a40013d50b032303a40013d58b02a302a40013d50b022302a40013d58b01a301a40013d50b012301a40013d58b00a300a4002300740113558d03a307a40013550d032307a40013558d02a306a40013550d022306a40013558d01a305a40013550d012305a40013558d00a304a4002304a40113d58a03a30ba40013d50a03230ba40013d58a02a30aa40013d50a02230aa40013d58a01a309a40013d50a012309a40013d58a00a308a40023085401c66a13d58c03a30fa40013d50c03230fa40013d58c02a30ea40013d50c02230ea40013d58c01a30da40013d50c01230da40013d58c00a30ca400230c940113050a16b305550192094e951396440097500000e780e0780529d29a23b48a1723b06a17231d2a21130da122930ba124cda76389a400814d19456397a4008144154929a0268919a0e5141949e2e09770ffffe7802023aa8a23380520231d05200355aa219349f9ffaa99239d3a2193155900d29503c6950183c6850103c7a50183c7b5012206558e4207e2075d8f598e83c6d50103c7c50183c7e50103c4f501a206d98ec2076204c18fdd8e8216558e233cc14603c6150183c6050103c7250183c735012206558e4207e2075d8f598e83c6550103c7450183c7650103c47501a206d98ec2076204c18fdd8e8216558e2338c14603c6950083c6850003c7a50083c7b5002206558e4207e2075d8f598e83c6d50003c7c50083c7e50003c4f500a206d98ec2076204c18fdd8e8216558e2334c14603c6150083c6050003c7250083c735002206558e4207e2075d8f598e83c6550003c7450083c7650083c57500a206d98ec207e205dd8dd58d8215d18d2330b146b14563e4b9006f30802dca8613041900018d630435016f30e02c5a8c6689930c0a161395460066950c65aee808612afc93155400d295139659005685368b97500000e780e01993154400e69513850a161396490097500000e7808018231d6a21033501468335814603360147833681472330a1362334b1362338c136233cd136528663930d0056860357a6219389140013945400329493974400ca8c628b637c370f2300740113d58b03a303a40013d50b032303a40013d58b02a302a40013d50b022302a40013d58b01a301a40013d50b012301a40013d58b00a300a4002304a40113558d03a307a40013550d032307a40013558d02a306a40013550d022306a40013558d01a305a40013550d012305a40013558d00a304a400a6652308b40013d58503a30ba40013d50503230ba40013d58502a30aa40013d50502230aa40013d58501a309a40013d505012309a40013d58500a308a400230c940113d58c03a30fa40013d50c03230fa40013d58c02a30ea40013d50c02230ea40013d58c01a30da40013d50c01230da40013d58c00a30ca40005aa139559003295b30d9740328913965d00a2853a8cbe8497500000e780e04713d58b03a303a40013d50b032303a40013d58b02a302a40013d50b022302a40013d58b01a301a40013d50b012301a40013d58b00a300a4002300740113558d03a307a40013550d032307a40013558d02a306a40013550d022306a40013558d01a305a40013550d012305a40013558d00a304a4002304a401a66513d58503a30ba40013d50503230ba40013d58502a30aa40013d50502230aa40013d58501a309a40013d505012309a40013d58500a308a4002308b40013d58c03a30fa40013d50c03230fa40013d58c02a30ea40013d50c02230ea40013d58c01a30da40013d50c01230da40013d58c00a30ca400230c940113050916b305950092094e9513964d0097500000e7804037a68762874a86c66de27486661b051700b305f60023b4d51623b06517231da62003358137833501370336813683360136233ca1782338b1782334c1782330d178233ca15a2338b15a2334c15a2330d15a03350a216309052c8149d687268c6e8d03598a218335815b0336015b8336815a0337015a233cb1782338c1782334d1782a8a2330e178835ba5212d4563ebab32cee4054b91491545bee0636fa9006309a900014b19456317a9000149954929a0ca8919a0651999499770ffffe780e0dbaa8a23380520231d05200355aa2113c4f9ffb30ca400239d9a2193955900d29503c6950183c6850103c7a50183c7b5012206558e4207e2075d8f598e83c6d50103c7c50183c7e50183c4f501a206d98ec207e204c58fdd8e8216558e233cc14603c6150183c6050103c7250183c735012206558e4207e2075d8f598e83c6550103c7450183c7650183c47501a206d98ec207e204c58fdd8e8216558e2338c14603c6950083c6850003c7a50083c7b5002206558e4207e2075d8f598e83c6d50003c7c50083c7e50083c4f500a206d98ec207e204c58fdd8e8216558e2334c14603c6150083c6050003c7250083c735002206558e4207e2075d8f598e83c6550003c7450083c7650083c57500a206d98ec207e205dd8dd58d8215d18d2330b146b14563e4bc006f20505f93841900058d630495016f20d05e13040a161395490022950c65aee8833d050093955400d29513965c00568597500000e78080d093954400a29513850a1613964c0097500000e78020cf231d3a21033501462330a13603358146833501470336814783dcaa212334a1362338b136233cc13613851c00b14563e4bc006f20704c33863b416304a6006f209057a66985098e04d2949385042213840a220e06228597500000e78040c9014593153500a2958c6133369501239ca5203295b3b6ac0093c61600758e23b8552165f2033581378335013703368136833601362334a1662330b166233cc1642338d1645285866763130b00568513060178ca85e2866a879770ffffe78040bb033501658335816503360166833681662330a15a2334b15a2338c15a233cd15a03350a21d687ee846e8cc66d6e8de31005d411a081494a6419e06f2090516a699770ffffe78040b423380520231d052023308522930519002338a420231c04202ae92eed130da122930ba124630439016f20d04e8355a52129466374b6006f20904e1b861500231dc520139655008336015b2a960337015a8337815b14ea8336815a18e21cee1307052214e6139645002a96233096162334b6178505139635003a962330560123b8aa20239cba2039a8130601785285ca85e2866a879770ffffe78000ad130da122930ba124854d930a40088a7585052ef1327592757266d2662aeb2ee732e3b6fe280b0c1a1306200497500000e780c0b1034481177d461305111e9305911797500000e78060b0814c81491375e40f2300a11e05447e75de75233ca1203e751e762338b120667c2334a120a2e42330c120230031230949630a0c2a0a68e28283d8625b01451387825b93975800b30517013383f5001386725d63036706aa830345070293f5f90fb3b4a5002d8d3335a000b3059040c98d95e501541305f121b28421c88345050083c70400b3b6f500bd8db335b000b306d040d58dfd147d150504e5d1138513001307170213061602e385b5fb13f5f50f09cd631608003da4c683630508228e039e9283b282727d1885bf33855303169583458500930485006387052003c5b40183c5a40103c6c40183c6d40122054d8d4206e206558e518d83c5f40103c6e40183c6040203c71402a205d18dc2066207d98ed58d82154d8d233ca17803c5340183c5240103c6440183c6540122054d8d4206e206558e518d83c5740103c6640183c6840103c79401a205d18dc2066207d98ed58d82154d8d2338a17803c5b40083c5a40003c6c40083c6d40022054d8d4206e206558e518d83c5f40003c6e40083c6040103c71401a205d18dc2066207d98ed58d82154d8d2334a17803c5340083c5240003c6440083c6540022054d8d4206e206558e518d83c5740003c6640083c6840003c79400a205d18dc2066207d98ed58d82154d8d2330a17803c5b40383c5a40303c6c40383c6d40322054d8d4206e206558e518d83c5f40303c6e40383c6040403c71404a205d18dc2066207d98ed58d82154d8d2334a16603c5340383c5240303c6440383c6540322054d8d4206e206558e518d83c5740303c6640383c6840303c79403a205d18dc2066207d98ed58d82154d8d2330a16603c5b40283c5a40203c6c40283c6d40222054d8d4206e206558e518d83c5f40203c6e40283c6040303c71403a205d18dc2066207d98ed58d82154d8d233ca16403c5340283c5240203c6440283c6540222054d8d4206e206558e518d83c5740203c6640283c6840203c79402a205d18dc2066207d98ed58d82154d8d2338a16403c41400054931a8c9a403c4140093852400130501787d4697500000e780a080014903c524046306052003c5d40583c5c40503c6e40583c6f40522054d8d4206e206558e518d83c5140603c6040683c6240603c73406a205d18dc2066207d98ed58d82154d8d233ca14603c5540583c5440503c6640583c6740522054d8d4206e206558e518d83c5940503c6840583c6a40503c7b405a205d18dc2066207d98ed58d82154d8d2338a14603c5d40483c5c40403c6e40483c6f40422054d8d4206e206558e518d83c5140503c6040583c6240503c73405a205d18dc2066207d98ed58d82154d8d2334a14603c5540483c5440403c6640483c6740422054d8d4206e206558e518d83c5940403c6840483c6a40403c7b404a205d18dc2066207d98ed58d82154d8d2330a14603c5d40783c5c40703c6e40783c6f40722054d8d4206e206558e518d83c5140803c6040883c6240803c73408a205d18dc2066207d98ed58d82154d8d233ca13603c5540783c5440703c6640783c6740722054d8d4206e206558e518d83c5940703c6840783c6a40703c7b407a205d18dc2066207d98ed58d82154d8d2338a13603c5d40683c5c40603c6e40683c6f40622054d8d4206e206558e518d83c5140703c6040783c6240703c73407a205d18dc2066207d98ed58d82154d8d2334a13603c5540683c5440603c6640683c6740622054d8d4206e206558e518d83c5940603c6840683c6a40603c7b406a205d18dc2066207d98ed58d82154d8d2330a13683ca3404054b29a883ca340493854404130501467d4697400000e780205e014b03358179833501790336817883360178233ca15a2338b15a2334c15a2330d15a033501658335816503360166833681662338a126233cb1262330c1282334d128033501468335814603360147833681472334a1222338b122233cc1222330d124033581378335013703368136833601362338a1762334b1762330c176233cd1740335815b8335015b0336815a8336015a233ca1782338b1782334c1782330d178033501278335812703360128833681282338a164233cb1642330c1662334d166033581228335012303368123833601242338a172233cb1722330c1742334d174033501778335817603360176833681752330a172233cb1702338c1702334d170139a8903cee893f9790009456312a9041355ba03ac1a2e9503450500335535010589930a4008630a052c1305015a7d46814597400000e780803d88162c0b1306200497400000e7806049014a0149f1a1a28d230081469305017813060002130401781305114697400000e78020479305016513060002930401651305114897400000e780a045a300614b2301514b93050173130600021305314a97400000e780e04393058170130600021305314c97400000e780a0421355ba036e8aac1a2e95034505003355350105892c0b19e903498119034a91191304a1199304a11b9305114a03459401034684018346a4010347b4012205518dc2066207d98e558d0346d4018346c4010347e4018347f4012206558e4207e2075d8f598e0216518d233ca15a034514010346040183462401034734012205518dc2066207d98e558d034654018346440103476401834774012206558e4207e2075d8f598e0216518d2338a15a03459400034684008346a4000347b4002205518dc2066207d98e558d0346d4008346c4000347e4008347f4002206558e4207e2075d8f598e0216518d2334a15a034514000346040083462400034734002205518dc2066207d98e558d034654008346440003476400834774002206558e4207e2075d8f598e0216518d2330a15a03c5940003c6840083c6a40003c7b4002205518dc2066207d98e558d03c6d40083c6c40003c7e40083c7f4002206558e4207e2075d8f598e0216518d2330a17603c5140103c6040183c6240103c734012205518dc2066207d98e558d03c6540183c6440103c7640183c774012206558e4207e2075d8f598e0216518d2334a17603c5940103c6840183c6a40103c7b4012205518dc2066207d98e558d03c6d40183c6c40103c7e40183c7f4012206558e4207e2075d8f598e0216518d2338a17603c5140003c6040083c6240003c734002205518dc2066207d98e558d03c6540083c6440003c7640083c774002206558e4207e2075d8f598e0216518d233ca17488161306200497400000e780001f930a4008c669854d15a4034981199307a11903c5170083c5070003c6270083c6370022054d8d4206e206558e518d83c5570003c6470083c6670003c77700a205d18dc2066207d98ed58d82154d8d2330a15a03c5970083c5870003c6a70083c6b70022054d8d4206e206558e518d83c5d70003c6c70083c6e70003c7f700a205d18dc2066207d98ed58d82154d8d2334a15a03c5170183c5070103c6270183c6370122054d8d4206e206558e518d83c5570103c6470183c6670103c77701a205d18dc2066207d98ed58d82154d8d2338a15a03c5970183c5870103c6a70183c6b70122054d8d4206e206558e518d83c5d70103c6c70183c6e70103c7f701a205d18dc2066207d98ed58d82154d8d233ca15a9307a11b03c5970083c5870003c6a70083c6b70022054d8d4206e206558e518d83c5d70003c6c70083c6e70003c7f700a205d18dc2066207d98ed58d82154d8d2330a17603c5170183c5070103c6270183c6370122054d8d4206e206558e518d83c5570103c6470183c6670103c77701a205d18dc2066207d98ed58d82154d8d2334a17603c5970183c5870103c6a70183c6b70122054d8d4206e206558e518d83c5d70103c6c70183c6e70103c7f701a205d18dc2066207d98ed58d82154d8d2338a17603c5170083c5070003c6270083c6370022054d8d4206e20683c55700558e518d03c64700a20583c6670003c77700d18d034a9119c2066207d98ed58d82154d8d233ca174881613061002814597400000e78080efc66923042123a30441239305015a130600026a8597400000e780a0fa93058175130600025e8597400000e78080f9881c8c161306200497400000e78080f8630c0920281d0c041306100297400000e78040f703451d0083450d0003462d0083463d0022054d8d4206e206558e518d83455d0003464d0083466d0003477d00a205d18dc2066207d98ed58d82154d8d2330a17803459d0083458d000346ad008346bd0022054d8d4206e206558e518d8345dd000346cd008346ed000347fd00a205d18dc2066207d98ed58d82154d8d2334a17803451d0183450d0103462d0183463d0122054d8d4206e206558e518d83455d0103464d0183466d0103477d01a205d18dc2066207d98ed58d82154d8d2338a17803459d0183458d010346ad018346bd0122054d8d4206e206558e518d8345dd010346cd018346ed010347fd01a205d18dc2066207d98ed58d82154d8d233ca17803c59b0083c58b0003c6ab0083c6bb0022054d8d4206e206558e518d83c5db0003c6cb0083c6eb0003c7fb00a205d18dc2066207d98ed58d82154d8d233ca16403c51b0183c50b0103c62b0183c63b0122054d8d4206e206558e518d83c55b0103c64b0183c66b0103c77b01a205d18dc2066207d98ed58d82154d8d2330a16603c59b0183c58b0103c6ab0183c6bb0122054d8d4206e206558e518d83c5db0103c6cb0183c6eb0103c7fb01a205d18dc2066207d98ed58d82154d8d2334a16603c51b0083c50b0003c62b0083c63b0022054d8d4206e206558e518d83c55b0003c64b0083c66b0003c77b00a205d18dc2066207d98ed58d82154d8d2338a164054b95a01795feff9305c542130600021305912297400000e78000188345012701254d8d05e11795feff9305a540130600021305112797400000e780e01501256309055c281d0c041306100297400000e78000d2130501787d46ea8597400000e78000d1014be6e003450127630a05209307212703c5970183c5870103c6a70183c6b70122054d8d4206e206558e518d83c5d70103c6c70183c6e70103c7f701a205d18dc2066207d98ed58d82154d8d233ca14603c5170183c5070103c6270183c6370122054d8d4206e206558e518d83c5570103c6470183c6670103c77701a205d18dc2066207d98ed58d82154d8d2338a14603c5970083c5870003c6a70083c6b70022054d8d4206e206558e518d83c5d70003c6c70083c6e70003c7f700a205d18dc2066207d98ed58d82154d8d2334a14603c5170083c5070003c6270083c6370022054d8d4206e206558e518d83c5570003c6470083c6670003c77700a205d18dc2066207d98ed58d82154d8d2330a1469307212903c5970083c5870003c6a70083c6b70022054d8d4206e206558e518d83c5d70003c6c70083c6e70003c7f700a205d18dc2066207d98ed58d82154d8d2334a13603c5170183c5070103c6270183c6370122054d8d4206e206558e518d83c5570103c6470183c6670103c77701a205d18dc2066207d98ed58d82154d8d2338a13603c5970183c5870103c6a70183c6b70122054d8d4206e206558e518d83c5d70103c6c70183c6e70103c7f701a205d18dc2066207d98ed58d82154d8d233ca13603c5170083c5070003c6270083c6370022054d8d4206e206558e518d83c5570003c6470083c6670003c77700a205d18dc2066207d98ed58d8215034911274d8d2330a136854c29a803491127130501467d469305212797400000e780e0ad814c03358179833501790336817883360178233ca1342338b1342334c1342330d134033501658335816503360166833681662330a1322334b1322338c132233cd132033501468335814603360147833681472330a1302334b1302338c130233cd13003358137833501370336813683360136233ca12e2338b12e2334c12e2330d12e63030c028a642c1d62859770ffffe780c0ba2e8471c5638604120e046294033c8472fd14cdb7900508622330a15608660c6a030686018334812b2334a1562338b156230cc1569770ffffe780809f833501562a84233c955a033581562330b45c83350157233004002334a45c030581572338b45c8544231b945a230ca45c23046401a30444011305a4008c061306000297400000e780409c1305a4020c161306000297400000e780209b23059405a30524051305c4040c061306000297400000e78080991305c4068c151306000297400000e7806098a2fc02e1866c6f001002330554032a9c23046c01a3044c011305ac008c061306000297400000e780c0951305ac020c161306000297400000e780a09423059c05a3052c051305cc040c061306000297400000e78000931305cc068c151306000297400000e780e091866c7daf4afc940588628c66906a83c686012330a1562334b1562338c156230cd156230cd1582338c1582334b1582330a15883596c5b0339812b2d4563f9a906da8dd28b13058c5b130b140093145400b3058500ae94330a540363fc69072380240113558903a383a400135509032383a40013558902a382a400135509022382a40013558901a381a400135509012381a40013558900a380a4001385840093050158654697400000e78020876da0930b4008054d914a154552f85af46369a4126303a412014d19456311a4120144954a39aa93155b005a952e9533848940131654002296a68597400000e780e0c713558903a383a400135509032383a40013558902a382a400135509022382a40013558901a381a400135509012381a40013558900a380a400238024011385840093050158654697300000e780207e13058c00b305450133065b0332953306540397400000e78060c18529629a2304ba01a3047a011305aa008c061306000297300000e780a07a1305aa020c161306000297300000e780807923059a056275a305aa041305ca040c061306000297300000e780c0771305ca068c151306000297300000e780a076231b3c5b854d6da463020c600a653384ad400c0462859770ffffe780e08a630f05586305b45f8e05e29503bc85720504cdb7a28a19a06514994a9760ffffe78020712a8b23300500231b055a83596c5b93c4faffce94231b955a930d8c5b93955a0033855d01aa95130501651306100297300000e780206f130a8c0033857a035295834b050093051500130501781306300897300000e780006d314563e4a4006f10a06c66f0ea8c138d1a003385a941630495006f10e07213058b5b93155d00ea9dee9513965400269697300000e780806913064008b305cd02d29513058b003386c40297300000e780e067231b5c5b1305015a930501651306100297300000e780606613050146930501781306300897300000e7802065628d63930c005a8d83596d5b13058d5b930d140093145400b3058500ae94930a4008330a540363fab9052380240113558903a383a400135509032383a40013558902a382a400135509022382a40013558901a381a400135509012381a40013558900a380a4001385840093050158654697300000e780a05d59a093955d006e952e9533848940131654002296a68597400000e780a0a013558903a383a400135509032383a40013558902a382a400135509022382a40013558901a381a400135509012381a40013558900a380a400238024011385840093050158654697300000e780e05613058d00b305450133865d0332953306540397400000e780209a854d027485296a9a22752304aa004275a304aa001305aa008c061306000297300000e780e0521305aa020c161306000297300000e780c05123058a046275a305aa041305ca040c061306000297300000e78000501305ca068c151306000297300000e780e04e231b3d5b130581759305015a1306100297300000e780604d8816930501461306600897300000e780404c130da12209456397ab00930ba124866cc669b9a613058162930581751306100297300000e780c0491305015a8c161306300897300000e780a04803350c00c669014a630705225a84835c4c5b2a8c13058170930581621306100297300000e7802046230071479305015a130630081305114697300000e780a044630400006f10804783596c5b2d4563eba92a52fc854d114a154522f8930b400863efac006389ac00814d19456397ac00814c154a29a0668a19a0e51c194a9760ffffe78060412a8b23300500231b055a03596c5b9344faffca94231b955a930a8c5b93155a0033854a01aa95130581751306100297300000e780e03c13048c0033057a032295034d05009305150088161306300897300000e780e03a314563e4a4006f10803aee8b930d1a003305b941630495006f10603d13058b5b93955d00ee9ad69513965400269697300000e7808037930a4008b3855d03a29513058b003386540397300000e780e035231b4c5b13050173930581751306100297300000e7806034130501788c161306300897300000e780403303546b5b13051400b1456364b4006f10c032338649416304a6006f104036627a050a8e0de29d93858d7293048b720e06268597300000e780a02f014593153500a6958c6133368500239aa55a3295b336a40093c61600758e23b0650165f21305016e930501731306100297300000e780202c13050165930501781306300897300000e780e02a6285854dc66963930b005a851306817093060146e68542779760ffffe780802c0945630fad10ea8b130581629305016e1306100297300000e78020271305015a930501651306300897300000e780e02503350c005a84e31e05dce67499e06f10e02d0a699760ffffe78040252a8423300500231b055a233495721305190080e0239a045aa2fc2ae1130da122866c630449016f10402b8354645b2945637495006f10402b130984721b851400231ba45a13955400b30594002e951305855b930581621306100297300000e780001e3385540322952304750125059305015a1306300897300000e780401c8504139534004a952330650123308b00231a9b5aa1a02300015a631eb40923308137233401362338b136130501468c161306015a9760ffffe780203559aa13068170930601466285e68522879760ffffe780a01ac669130da122866c930ba124aa64850426e57e75de753e769e762aeb2ee732e3b6fe280b90133414981cce8597a0ffffe780009d13f51c00631e0516a66413f5f40f130515f0933c1500138414008813ac1a26869750ffffe780c0e3a6896fe0afe18e05e29503b5857219c8b30580400356655b0e06329503358572fd15edf98355655bfd152338a164233c01642330b16613050146930501651306015a9760ffffe780402913050178930501461306500a97300000e780600b03358150033a81518355655b03340151aa84636fba00046191c8035a455b83d5645b05042685e378bafe19a0228a2a8413155a00b38544012e959309855b33055a03269513098500881613061002ce8597300000e780e00593050178130610024e8597300000e780c0041306400813051138ca8597300000e780a003130640084a859305117a97300000e780800209cc0e0ad29483b404737d14c66919c483b484727d146dfc11a0c669130501468c161306500a97300000e780a0ff23349150233801502a658345015a7d152ae5e38505e8667519e16f10200c8a6599e16f10400c03368572b2fcfd152ee12330060097f0feffe78000ad85b5a8082c0b97a0ffffe78000a16fd00ff92689aa84033a8148833a014813155900229583459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18d233cb13683451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2338b13683459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2334b13683451500034605008346250003473500a205d18dc20662070346550083474500d98ed58d22065d8e834665000347750093174900b309f400c2066207d98e558e0216d18d2330b136930501781306000297300000e78020e803b5891683b5091623b0591723b4491791cc0e094a9403348422fd14930a400881c803340422fd14edfc19a0930a400803368137833601370337813683370136233cc1462338d1462334e1462330f1462330b1482334a14823388148233c01480a758345015a7d152af199e16fe0afad4a65e30d0570ea65e38f05700336052232e9fd152eed2338062097f0feffe78020906fe04fabe6650676a6762eef467732f336f7e6753afb2a660a643339b000b3062041b3f9c600638d09063336200193361500758e11ca054909c483b585727d146dfc014a2e8521a02e8ae30a09668355655b6362b4020461e381045a0354455b050a97f0feffe780808983d5645b2685e373b4fe26858145fd190504e3050afa0e042295033585729304faff81450144d9d803358572fd14edfc8145014461b7630a090219e52e8509c4033585727d146dfc0c6191c92e8497f0feffe78020840c602285edf911a02a84228597f0feffe780e082ca6501450a766a6a3339b000b3062041b3f9c600638e09063336200193361500758e01ce054963070a0083b505227d1ae31d0afe81442e8521a0ae84e30c095a8355a5216363ba0203340521e306044e035a8521850497e0feffe780007d8355a4212285e372bafe22858145fd19050ad5d00e0a529503350522fd148145014ad1d803350522fd14edfc8145014a59b7630e090209e92e8563070a00033505227d1ae31d0afe8335052199c92e8497e0feffe7808077833504212285e5f911a02a84228597e0feffe780207613050004854597e0feffe780c074e3040558aa8dc26703c5970183c5870103c6a70183c6b70122054d8d4206e206558e518d83c5d70103c6c70183c6e70103c7f701a205d18dc2066207d98ed58d82154d8d233ca14603c5170183c5070103c6270183c6370122054d8d4206e206558e518d83c5570103c6470183c6670103c77701a205d18dc2066207d98ed58d82154d8d2338a14603c5970083c5870003c6a70083c6b70022054d8d4206e206558e518d83c5d70003c6c70083c6e70003c7f700a205d18dc2066207d98ed58d82154d8d2334a14603c5170083c5070003c6270083c6370022054d8d4206e206558e518d83c5570003c6470083c6670003c77700a205d18dc2066207d98ed58d82154d8d2330a146130501482c0b1306000297300000e78080b293050146130600046e8597300000e78060b185458546854c6e8501469770ffffe780409d6265033c050109452afa02fe82e2e3090c280949014b014482e46265033a05001785feff1305e598aae893044006130d00108949b3058a0003c50500130685fba546e3eec62a0e06c66636961062930a14000286e36f2b23d27933059b024e950344e5fb130940068944e307943e1306c5f9835bc5f90355c6018355a6018356e6010357060242054d8d82164217d98e558d2334a1280355460183552601835666010357860142054d8d82164217d98e558d2330a1280355c6008355a60042058356e600035706014d8d9305360282164217d98e558d233ca126035546008356260003576600035686004205558d02174216598e518d2338a126130610041305117897300000e780a09f23008178791bdae233052b034e95034425020949e3029434835405008355c5010356a5018356e50103570502c205d18d82164217d98ed58daee183554501035625018356650103578501c205d18d82164217d98ed58d2efd8355c5000356a500c2058356e500035705014d8e9305350282164217d98e558e32f9035645008356250003576500035585004206558e02174215598d518d2af5130610041305113697300000e780209533c574011335150093b50b106d8d23008136e307050ca8082c115e869740ffffe78060651305015a8c1c5e869740ffffe7806064a8089305015a1306000297300000e78040d30125e31c050813958b036d912c112e950345050093f57b003355b5000589630d056c13050146b008930601789816d9ad2665e314050626651a056e9583459501034685018346a5010347b501a205d18dc2066207d98ed58d0346d5018346c5010347e5018347f5012206558e4207e2075d8f598e0216d18d233cb14683451501034605018346250103473501a205d18dc2066207d98ed58d034655018346450103476501834775012206558e4207e2075d8f598e0216d18d2338b14683459500034685008346a5000347b500a205d18dc2066207d98ed58d0346d5008346c5000347e5008347f5002206558e4207e2075d8f598e0216d18d2334b14683451500034605008346250003473500a205d18dc2066207d98ed58d034655008346450003476500834775002206558e4207e2075d8f598e0216d18d2330b14683459503034685038346a5030347b503a205d18dc2066207d98ed58d0346d5038346c5030347e5038347f5032206558e4207e2075d8f598e0216d18d233cb13683451503034605038346250303473503a205d18dc2066207d98ed58d034655038346450303476503834775032206558e4207e2075d8f598e0216d18d2338b13683459502034685028346a5020347b502a205d18dc2066207d98ed58d0346d5028346c5020347e5028347f5022206558e4207e2075d8f598e0216d18d2334b13683451502034605028346250203473502a205d18dc2066207d98ed58d034655028346450203476502034575022206558e42076205598df276518d02154d8d2330a1366319db00081ada859790ffffe78040ec166bd27933059b023384a9002310040013052400930501461306000297200000e780a06923010402130534028c161306000297200000e7804068050bdae226650505aae4f9a133356001b3b58a016d8d630e055ed29a83ca0a0063940a00930a00107d1bdae233059b024e9583442502638b247b835c05008355c5010356a5018356e50103570502c205d18d82164217d98ed58d233cb13683554501035625018356650103578501c205d18d82164217d98ed58d2338b1368355c5000356a500c2058356e500035705014d8e9305350282164217d98e558e2334c136035645008356250003576500035585004206558e02174215598d518d2330a136130501461306100497200000e780205b03358137833501370336813683360136aaf8aef4b2f0b6ec2300917893050146130610041305117897200000e780205863f7ac514675a6750676e666233ca15a2338b15a2334c15a2330d15a63820a2c8144b38b9c0013950b0341916371a54f1305015aac085e869740ffffe780a02613958b036d91ac082e950345050093f57b003355b500058915c11305014613061002814597200000e780804488161306015a93060146130701780da01305014613061002814597200000e780604288161306015a9306017813070146de859790ffffe78000d78504130501788c161306200497200000e780804c139504034191e36155f739ac63050b44930b140263e48b50636f7c43637f746133855b4193050002631eb55cb3055a01130600021305117897200000e78080487d1bdae2d2792300017833059b024e958344250289456392b408dda3630d0b3e930b240463e18b4c63677c3f63f38a4d130524026360ac4c63e2ab5c130940063386ab4093060002631ed656d29a83c40a0013842500b305aa00130600021305217a97200000e780e0411306000213052178a28597200000e780c0407d1bdae2d279a30091782300917933052b034e95834425028945638ab456035405008355c5010356a5018356e50103570502c205d18d82164217d98ed58daef883554501035625018356650103578501c205d18d82164217d98ed58daef48355c5000356a500c2058356e500035705014d8e9305350282164217d98e558eb2f0035645008356250003576500035585004206558e02174215598d518daaec130610041305113697200000e780e035230091366374a42f1305015aac0822869740ffffe780e006131584036d91ac082e9503450500937574003355b500058909c9130501461306015a93060178981601a8130501461306015a941613070178a2859790ffffe78080b9930440067275631cab000949081ada859790ffffe78020af166bd27911a00949050433059b02b384a90023908400138524009305015a1306000297200000e780202c1385240293044006930501461306200497200000e780a02a050bdae2de8ae5a8e68b0335015a8335815a0336015b8336815b2330a1362334b1362338c136233cd13613050146930501781306200497200000e780c0267275631aab00081ada859790ffffe78000a6166bd279854c93044006930a2400850b33059b023384a90023107401130524008c161306000297200000e780c02213052402930501461306200497200000e7808021166b9da013050146b008941613070178de859790ffffe78020a9930440067275631aab00081ada859790ffffe780e09e166bd279850b33059b023384a9002310740113052400ac081306000297200000e780401c13052402930501461306200497200000e780001b050bdae2568463ed8aed05456319ab1252740355040013450510a66593c515004d8d631e051093052402130511659790ffffe780a0bd727511c5228597e0feffe780e0c76e8597e0feffe78040c703156165831541650356216583061165231aa172c205d18d033581662328b1728305016703348165233ca174833401662300b1762304d1221305912293050173194697200000e780801113558403230ba12213550403a30aa12213558402230aa12213550402a309a122135584012309a12213550401a308a122135584002308a122a307812213d58403230fa12213d50403a30ea12213d58402230ea12213d50402a30da12213d58401230da12213d50401a30ca12213d58400230ca122a30b91221305f12393058175254697200000e780e008281413060002a26597200000e780604a814c01251334150005a0854c727511c5527597e0feffe78060b76e8597e0feffe780c0b613044002e265886511c5886197e0feffe78080b56685a2850d618330817e0334017e8334817d0339017d8339817c033a017c833a817b033b017b833b817a033c017a833c8179033d0179833d81781301017f8280a308a16441bfad452685ada0b1459da097e0feffe78000b01775feff1305a56c09a897e0feffe780e0ae1775feff1305856b9305b00291a81785feff130515839305500399a01775feff1305b57f25a81775feff1305157f3da01775feff1305656b29a01775feff1305c56af14531a85685e2859730ffffe78040f500001775feff1305357c930580029720ffffe780a06900001775feff1305e56459bf1775feff1305257593050003c5b71775feff1305655f93050002c9bfad4566855dbf1775feff130515787dbf1775feff1305757755bf1775feff1305e56099bf1775feff13054560b1b71775feff1305a55f89b71775feff1305e5729305100271b7ad454e8585bf1775feff1305b573a5bf1775feff1305255d29bf1775feff13056570e1bf1775feff1305e55b19b71775feff1305256c85bf1775feff1305a55695bf13050002930500022db71305000497e0feffe780809d00001775feff13058558c1bd1775feff1305e557d9b51775feff1305455775bd5685de85e5bd1775feff1305455675b51775feff1305a5554db5034715008347050022075d8f83472500c207d98f0347350062075d8f834745008217d98f0347550022175d8f8347650003457500c217d98f62155d8d82802e869737000083b7675c814582870971a2faa6f6caf286feceeed2ead6e6dae25efe62fa66f66af26eee2ae4ae8401441309000833858400eff0bff8930704018a9788e32104e31724ffa265130600040809ef10d05d4a754a6fc2679782feff83b242942a9f3e9fa267e269ea78b4639787feff83b78795ea6eb346df00bd8e939706028192dd8eb692334555009357850122155d8d4e9f2a9fb346df0093d70601c216dd8eb69233c5a200931715007d915d8d8277c69e978ffeff83bf0f90be9ea2670e660a7eb8679787feff83b7678ec27b33c7ee003d8f9317070201935d8fba9fb3c8f80193d78801a218b3e8f800a277329e5e9ebe9ec69e33c7ee009357070142175d8fba9fb3c81f019397180093d8f803b3e8f800a2679785feff83b5c58b978cfeff83bc4c88bc6b2e682a73b347fe00ad8f939507028193cd8fbe9c334696019355860122164d8ee275066442932e9e329eb347fe0093d50701c217cd8fbe9c33c6cc00931516007d924d8ea26522939783feff83b3a384ac6d178dfeff033d0d85a664b345b300b3c57500939305028191b3e575002e9d3348a80193538801221833687800269342934669b345b30093d30501c215b3e575002e9d4a9f33480d01469f93131800b345bf001358f80333687800939305028191b3e57500666bae9cb3c81c0193d38801a218b3e878005a9f469f067ab345bf0093d30501c215b3e57500ae9cd29eb3c81c01b29e93931800b3c6de0093d8f803b3e87800939306028192b3e67600a674369d3346cd0093538601221633667600a69eb29eb3c6de0093d30601c216b3e67600369d3346cd00931316007d9233667600c673e67a0a6c1e9e429e3347ee00931407020193458fba9233c8020193548801221833689800569e429e3347ee00935407014217458fba92629333c802012a9393141800b347f3001358f80333689800939407028193c58fbe9f33c5af00935485012215458daa64629fde9e26932a93b347f30093dd0701c217b3e7b701be9f33c5af00931d15007d913365b5012a9fb346df00939d06028192b3e6b601b69233c5a200935d850122153365b501529f2a9fb346df0093dd0601c216b3e6b601b69233c5a200c69e931d150033c7ee007d913365b501931d070201933367b701ba9fb3c81f0193dd8801a218b3e8b801ca9ec69e33c7ee00935d070142173367b701ba9f5a9eb3c81f01329e939d1800b347fe0093d8f803b3e8b801939d07028193b3e7b701be9c33c6cc00935d860122163366b601269e329eb347fe0093dd0701c217b3e7b701be9c569333c6cc004293931d1600b345b3007d923366b601939d05028191b3e5b5012e9d33480d01935d880122183368b80122934293b345b30093dd0501c215b3e5b5012e9d4e9f33480d01469f931d1800b345bf001358f8033368b801939d05028191b3e5b501ae9cb3c81c0193dd8801a218b3e8b8011e9f469fb345bf0093dd0501c215b3e5b501ae9cb3c81c01939d180093d8f803b3e8b801c26dee9eb29eb3c6de00939d06028192b3e6b601369d3346cd00935d860122163366b601827dee9eb29eb3c6de0093dd0601c216b3e6b601369d3346cd00931d16007d923366b601a67d9e9ec69e6e9e429e3347ee00931d070201933367b701ba9233c80201935d880122183368b801a66d6e9e429e3347ee00935d070142173367b701ba9233c80201931d18001358f8033368b801e27d33c7ee006e932a93b347f300939d07028193b3e7b701be9f33c5af00935d850122153365b501a27d6e932a93b347f30093dd0701c217b3e7b701be9f33c5af00931d15007d913365b501a67d269342936e9f2a9fb346df00939d06028192b3e6b601b69233c5a200935d850122153365b5014a9f2a9fb346df0093dd0601c216b3e6b601b69233c5a200931d15007d913365b501931d070201933367b701ba9fb3c81f0193dd8801a218b3e8b801c26db345b3005693ee9ec69e33c7ee00935d070142173367b701ba9fb3c81f01939d180093d8f803b3e8b801e27d529f469f6e9e329eb347fe00939d07028193b3e7b701be9c33c6cc00935d860122163366b601827d6e9e329eb347fe0093dd0701c217b3e7b701be9c33c6cc00931d16007d923366b601939d05028191b3e5b5012e9d33480d01935d880122183368b8014293b345b30093dd0501c215b3e5b5012e9d33480d01931d1800b345bf001358f8033368b801939d05028191b3e5b501ae9cb3c81c0193dd8801a218b3e8b801629f469fb345bf0093dd0501c215b3e5b501ae9cb3c81c01939d180093d8f803b3e8b801a27d5a932a93ee9eb29eb3c6de00939d06028192b3e6b601369d3346cd00935d860122163366b601a29eb29eb3c6de0093dd0601c216b3e6b601369d3346cd00931d16007d923366b601a66db347f3005e936e9e429e3347ee00931d070201933367b701ba9233c80201935d880122183368b8014e9e429e3347ee00935d070142173367b701ba9233c80201931d18001358f8033368b801939d07028193b3e7b701be9f33c5af00935d850122153365b5012a93b347f30093dd0701c217b3e7b701be9f33c5af00931d15007d913365b501a66d569e329e6e9f2a9fb346df00939d06028192b3e6b601b69233c5a200935d850122153365b5015a9f2a9fb346df0093dd0601c216b3e6b601b69233c5a200931d15007d913365b501a27db347fe001e9eee9ec69e33c7ee00931d070201933367b701ba9fb3c81f0193dd8801a218b3e8b801ce9ec69e33c7ee00935d070142173367b701ba9fb3c81f01939d180093d8f803b3e8b801939d07028193b3e7b701be9c33c6cc00935d860122163366b601329eb347fe0093dd0701c217b3e7b701be9c33c6cc00931d16007d923366b601a67d5e9e6e934293b345b300939d05028191b3e5b5012e9d33480d01935d880122183368b80162934293b345b30093dd0501c215b3e5b5012e9d33480d01931d18001358f8033368b801827d429e3347ee006e9f469fb345bf00939d05028191b3e5b501ae9cb3c81c0193dd8801a218b3e8b801229f469fb345bf0093dd0501c215b3e5b501ae9cb3c81c01939d180093d8f803b3e8b801e27d26932a93ee9eb29eb3c6de00939d06028192b3e6b601369d3346cd00935d860122163366b601d29eb29eb3c6de0093dd0601c216b3e6b601369d3346cd00931d16007d923366b601931d070201933367b701ba9233c80201935d880122183368b801c26db347f3004a936e9e429e3347ee00935d070142173367b701ba9233c80201931d18001358f8033368b801939d07028193b3e7b701be9f33c5af00935d850122153365b5012a93b347f30093dd0701c217b3e7b701be9f33c5af00931d15007d913365b5015a9f2a9fb346df00939d06028192b3e6b601b69233c5a200935d850122153365b501c26d529342936e9f2a9fb346df0093dd0601c216b3e6b601b69233c5a200931d15007d913365b501e27db345b3002693ee9ec69e33c7ee00931d070201933367b701ba9fb3c81f0193dd8801a218b3e8b801a66d629fee9ec69e33c7ee00935d070142173367b701ba9fb3c81f01939d180093d8f803b3e8b801827d469f6e9e329eb347fe00939d07028193b3e7b701be9c33c6cc00935d860122163366b6015e9e329eb347fe0093dd0701c217b3e7b701be9c33c6cc00931d16007d923366b601939d05028191b3e5b5012e9d33480d01935d880122183368b8014293b345b30093dd0501c215b3e5b5012e9d33480d01931d1800b345bf001358f8033368b801939d05028191b3e5b501ae9cb3c81c0193dd8801a218b3e8b8014e9f469fb345bf0093dd0501c215b3e5b501ae9cb3c81c01939d180093d8f803b3e8b801a67d229e429eee9eb29eb3c6de00939d06028192b3e6b601369d3346cd00935d860122163366b6019e9eb29eb3c6de0093dd0601c216b3e6b601369d3346cd00931d16003347ee007d923366b601931d070201933367b701ba9233c80201935d880122183368b8014a9e429e3347ee00935d070142173367b701ba9233c80201931d18001358f8033368b801a27da29ec69e6e932a93b347f300939d07028193b3e7b701be9f33c5af00935d850122153365b50156932a93b347f30093dd0701c217b3e7b701be9f33c5af00931d15007d913365b501827d33c7ee00d29e6e9f2a9fb346df00939d06028192b3e6b601b69233c5a200935d850122153365b5011e9f2a9fb346df0093dd0601c216b3e6b601b69233c5a200931d15007d913365b501931d070201933367b701ba9fb3c81f0193dd8801a218b3e8b801c69e33c7ee00935d070142173367b701ba9fb3c81f01939d180093d8f803b3e8b801c26d4a9342936e9e329eb347fe00939d07028193b3e7b701be9c33c6cc00935d860122163366b601a67db345b3005e9f6e9e329eb347fe0093dd0701c217b3e7b701be9c33c6cc00931d16007d923366b601939d05028191b3e5b5012e9d33480d01935d880122183368b801a27d469f269e6e934293b345b30093dd0501c215b3e5b5012e9d33480d01931d1800b345bf001358f8033368b801939d05028191b3e5b501ae9cb3c81c0193dd8801a218b3e8b801569f469fb345bf0093dd0501c215b3e5b501ae9cb3c81c01939d180093d8f803b3e8b801a66d429e3347ee00ee9eb29eb3c6de00939d06028192b3e6b601369d3346cd00935d860122163366b601e27d629e4e93ee9eb29eb3c6de0093dd0601c216b3e6b601369d3346cd00931d16007d923366b601931d070201933367b701ba9233c80201935d880122183368b801429e3347ee00935d070142173367b701ba9233c802012a93931d1800b347f3001358f8033368b801939d07028193b3e7b701be9f33c5af00935d850122153365b5015a932a93b347f30093dd0701c217b3e7b701be9f33c5af00931d15007d913365b5011e9f2a9fb346df00939d06028192b3e6b601b69233c5a200935d850122153365b501e27dce9ec69e6e9f2a9fb346df0093dd0601c216b3e6b601b69233c5a200931d150033c7ee007d913365b501931d070201933367b701ba9fb3c81f0193dd8801a218b3e8b801a69ec69e33c7ee00935d070142173367b701ba9f629eb3c81f01329e939d1800b347fe0093d8f803b3e8b801939d07028193b3e7b701be9c33c6cc00935d860122163366b601569e329eb347fe0093dd0701c217b3e7b701be9c5e9333c6cc004293931d1600b345b3007d923366b601939d05028191b3e5b5012e9d33480d01935d880122183368b80152934293b345b30093dd0501c215b3e5b5012e9d33480d01931d18001358f8033368b801c26da29eb29e6e9f469fb345bf00939d05028191b3e5b501ae9cb3c81c0193dd8801a218b3e8b801a66db3c6de005a9e6e9f469fb345bf0093dd0501c215b3e5b501ae9cb3c81c01939d180093d8f803b3e8b801939d06028192b3e6b601369d3346cd00935d860122163366b601a27d429e3347ee00ee9eb29eb3c6de0093dd0601c216b3e6b601369d3346cd00931d16007d923366b601931d070201933367b701ba9233c80201935d880122183368b801827d4a932a936e9e429e3347ee00935d070142173367b701ba9233c80201931d1800b347f3001358f8033368b801939d07028193b3e7b701be9f33c5af00935d850122153365b501a67d569f1e9e6e932a93b347f30093dd0701c217b3e7b701be9f33c5af00931d15007d913365b5012a9fb34ddf0093960d0293dd0d02b3eddd00ee92b3c6a20013d58601a216c98e2675329eb347fe002a9f369fb34dbf0113d50d01c21db3edad00ee92b3c6d20013951600fd92c98e26654e9eaa9ec69e33c7ee00131507020193498fba9fb3c81f0113d58801a218b3e8a800e29ec69e33c7ee00135507014217498fba9fb3c81f011395180093d8f803b3e8a800139507028193c98fbe9c33c6cc00135586012216498e329eb347fe0013d50701c217c98fbe9c33c6cc00131516007d92498e2275a69eb29e2a934293b345b300139505028191c98d2e9d33480d011355880122183368a8005a934293b345b30013d50501c215c98d2e9d33480d01131518001358f8033368a8006275b3cdbe01de9e2a9f469fb345bf00139505028191c98dae9cb3c81c0113d58801a218b3e8a80042654a9e429e2a9f469fb345bf0013d50501c215c98dae9cb3c81c011395180093d8f803b3e8a80013950d0293dd0d02b3edad006e9d3346cd00135586012216498eb29eb3cdbe0113d50d01c21db3edad006e9d3346cd00131516003347ee007d92498e131507020193498fba9233c802011355880122183368a800229e429e3347ee00135507014217498fba9233c80201131518001358f8033368a8000275229fe29e2a933693b347f300139507028193c98fbe9fb3c6df0013d58601a216c98e52933693b347f30013d50701c217c98fbe9fb3c6df0013951600fd92c98e369fb34dbf0113950d0293dd0d02b3edad00ee92b3c6d20013d58601a216c98e269f369fb34dbf0113d50d01c21db3edad00ee92b3c6d200c69e1395160033c7ee00fd92c98e131507020193498fba9fb3c81f0113d58801a218b3e8a800da9ec69e33c7ee00135507014217498fba9fb3c81f011395180093d8f803b3e8a80026751e9f469f2a9e329eb347fe00139507028193c98fbe9c33c6cc00135586012216498e2275d69e2a9e329eb347fe0013d50701c217c98fbe9c33c6cc00131516007d92498e4265b29eb3cdbe012a934293b345b300139505028191c98d2e9d33480d011355880122183368a8004a934293b345b30013d50501c215c98d2e9d33480d0113151800b345bf001358f8033368a800139505028191c98dae9cb3c81c0113d58801a218b3e8a80002754e9e429e2a9f469fb345bf0013d50501c215c98dae9cb3c81c011395180093d8f803b3e8a80013950d0293dd0d02b3edad006e9d3346cd00135586012216498e26653347ee005e9eaa9eb29eb3cdbe0113d50d01c21db3edad006e9d3346cd00131516007d92498e131507020193498fba9233c802011355880122183368a800429e3347ee00135507014217498fba92529333c80201369313151800b347f3001358f8033368a800139507028193c98fbe9fb3c6df0013d58601a216c98e6275529fca9e2a933693b347f30013d50701c217c98fbe9fb3c6df0013951600fd92c98e369fb34dbf0113950d0293dd0d02b3edad00ee92b3c6d20013d58601a216c98e0275c69e33c7ee002a9f369fb34dbf0113d50d01c21db3edad00ee92b3c6d20013951600fd92c98e131507020193498fba9fb3c81f0113d58801a218b3e8a800de9ec69e33c7ee00135507014217498fba9fb3c81f011395180093d8f803b3e8a80026654e9342932a9e329eb347fe00139507028193c98fbe9c33c6cc00135586012216498e229e329eb347fe0013d50701c217c98fbe9c33c6cc0013151600b345b3007d92498e139505028191c98d2e9d33480d011355880122183368a8006275269f469f2a934293b345b30013d50501c215c98d2e9d33480d0113151800b345bf001358f8033368a800139505028191c98dae9cb3c81c0113d58801a218b3e8a8002675da9eb29e2a9f469fb345bf0013d50501c215c98dae9cb3c81c0113951800b3cdbe0193d8f803b3e8a80013950d0293dd0d02b3edad006e9d3346cd00135586012216498ee29eb29eb3cdbe0113d50d01c21db3edad006e9d3346cd00131516007d92498e2275569336932a9e429e3347ee00131507020193498fba9233c802011355880122183368a8001e9e429e3347ee00135507014217498fba9233c8020113151800b347f3001358f8033368a800139507028193c98fbe9fb3c6df0013d58601a216c98e42655e9e329e2a933693b347f30013d50701c217c98fbe9fb3c6df0013951600fd92c98e4265b347fe0022932a9f369fb34dbf0113950d0293dd0d02b3edad00ee92b3c6d20013d58601a216c98e4e9f369fb34dbf0113d50d01c21db3edad00ee92b3c6d20013951600fd92c98e02754293b345b300aa9ec69e33c7ee00131507020193498fba9fb3c81f0113d58801a218b3e8a80022754a9faa9ec69e33c7ee00135507014217498fba9fb3c81f011395180093d8f803b3e8a800139507028193c98fbe9c33c6cc00135586012216498e6275469fd29e2a9e329eb347fe0013d50701c217c98fbe9c33c6cc00131516007d92498e139505028191c98d2e9d33480d011355880122183368a8002665b29eb3cdbe012a934293b345b30013d50501c215c98d2e9d33480d0113151800b345bf001358f8033368a800139505028191c98dae9cb3c81c0113d58801a218b3e8a8005a9f469fb345bf0013d50501c215c98dae9cb3c81c011395180093d8f803b3e8a80013950d0293dd0d02b3edad006e9d3346cd00135586012216498e26751e9e429eaa9eb29eb3cdbe0113d50d01c21db3edad006e9d3346cd00131516003347ee007d92498e131507020193498fba9233c802011355880122183368a800569e429e3347ee00135507014217498fba92629333c80201369313151800b347f3001358f8033368a800139507028193c98fbe9fb3c6df0013d58601a216c98e26933693b347f30013d50701c217c98fbe9fb3c6df0013951600fd92c98e7a9c369cb34dbc0113950d0293dd0d02b3edad00ee92b3c6d20013d58601a216c98e629a369ab34dba0113d50d01c21db3edad00ee92f69bb3c6d200c69b1395160033c7eb00fd92c98e131507020193498fba9fb3c81f0113d58801a218b3e8a8005e9946993347e900135507014217498fba9f729bb3c81f01329b13951800b347fb0093d8f803b3e8a800139507028193c98fbe9c33c6cc00135586012216498eda94b294a58f13d50701c217c98fbe9c9a9a33c6cc00c29a13151600b3c5ba007d92498e139505028191c98d2e9d33480d011355880122183368a80056944294a18d13d50501c215c98d2e9dd29933480d01c69913151800b3c5b9001358f8033368a800139505028191c98dae9cb3c81c0113d58801a218b3e8a800ce93c6931ee9b3c3b30093d50301c213b3e3b3009e9ce6f1b3cc1c0193951c0093dcfc03b3e595012efdc2651ee6ca95b295b3cdb50113950d0293dd0d02b3edad006e9d3346cd00135586012216498e0275aa95b2952eedb3c5b50113d50501c215c98d2e9deaf5334dcd0013161d00135dfd033366a601b2e12676aef926964296318f1315070293550702c98dae9233c802011357880122183368e8002667329742973af12d8f135607014217518fba9296e9b3c20201bafd1397120093d2f20333675700bae5627722973697b98f9395070213d607024d8eb29fb3c6df0093d78601a216dd8ea277ba97b6973ef5b18f13d70701c217d98fbe9ffeedb3cfdf003ee293971f0093dfff03b3e7f7013ef9a26714091386070498638c62a107a1062d8f8c7e2d8f23bce7fee317f6fef6705674b6741679f669566ab66a166bf27b527cb27c127df26d19618280397156e4833a050e52e8130a000822f826f44af04eec06fc330a5a412a842e89b284930905066373ca0452862330050e33855901ef00a0323c603864938404f8938707083ce093b70708ba9752993ce4ce852285d694efe08fceb30a9900130a0008b3859a402e8963649a0268702686ca854e95ef00a02e7c70e2700279a6977cf04274a274e269426aa26a216182803c6038642285938707083ce093b70708ba973ce4efe0afc9938404f85dbf797122f04ae82a842e891306800b81451305050426ec4ee406f4ef00801c9767feff83b747e01ce09767feff83b727e11ce49767feff83b787df1ce89767feff83b767e11cec9767feff83b747e01cf09767feff83b727de1cf49767feff83b707e01cf89767feff83b7e7dd1cfc81449309000433059900efe0cfbc330794001c63a104a98f1ce3e39634ff83470900a270e2647cf402744269a269014545618280357122e926e54ae106ed2a84b2843689eff0fff4634805021306000881450a85ef0000124a86a6850a85ef00401e8a85228513060008eff0bfe7930500080a85efe00fbaea604a64aa640a6901450d61828009ca411106e4eff09fe5a260014541018280014582801d71a2e8a6e4cae02a84ae843289814513068003280086ec02e0ef00e00b7d55d5c47c747d556363f90a3c68c5e368703c603864aa973ce0b3b7a700ba973ce48347040f99c3fd573cecfd571309040613060008098e3ce881454a95ef00c007ca852285efe02fb28a87a286130604043e899862a106a10793558700a38cb7fe93550701238db7fe93558701a38db7fe93550702238eb7fe93558702238ce7fea38eb7fe935507036193238fb7fea38fe7fee390c6fc7074ca852685ef00a00e4a8593050004efe02fab0145e6604664a66406692561828071c693f7f50f2300f5003307c500a30ff7fe894663fcc60aa300f5002301f500230ff7fea30ef7fe994663f1c60aa301f500230ef7fea14663fac60893f5f50f9b9785003307a0400d8bad9f198e9b950701ad9f2a97719a1cc3b305c70023aef5fe63f5c6065cc31cc723aaf5fe23acf5fee14663fcc604137847005cc71ccb5ccb1ccf6108939807029396070293d8080223a2f5fe23a4f5fe23a6f5fe23a8f5fe33060641fd474297c69663f0c7020116937706fe93870702ba9714e314e714eb14ef13070702e31af7fe8280397122fc26f84af44ef052ec56e85ae45ee093f735006387074069c2aa8719a06303062a83c60500850513f735002380d7007d1685076df793f637003e87cdea3d48637dc804930806ff6378180133e8b700137878006304083093d84800138f1800120f2e9f2e87be86832e0700032e4700032387000328c70023a0d60123a2c60123a4660023a606014107c106e31eeffc85089208c695c6973d8a137886001377460093762600058a630c080083a8050003a84500a107a10523ac17ff23ae07ff11c798419107910523aee7fe6391061e09c603c705002380e7006274c27422798279626ac26a226b826b216182807d476379c70a094883c805009841638806290d486386061d9306c6fe03c3150003c8250093f306ff13843700938435009382330123801701a38067002381070113d94600ae92a687a28803a8170083a5570083a697001b53870103a7d7009b1f88001b9f85009b9e86001b5888019bd585019bd686011b1e87003363f3013368e801b3e5d501b3e6c60123a0680023a2080123a4b80023a6d800c107c108e39657fa9307190092073516b385f40033067640a29793780601137886009376460013772600058a6384080883cb050003cb150083ca250003ca350083c9450003c9550083c4650003c4750083c3850083c2950083cfa50003cfb50083cec50003ced50003c3e50083c8f50023807701a380670123815701a381470123823701a382270123839700a383870023847700a38457002385f701a385e7012386d701a386c70123876700a3871701c105c1076304080483c2050083cf150003cf250083ce350003ce450003c3550083c8650003c8750023805700a380f7012381e701a381d7012382c701a382670023831701a3830701a105a1079dc203c3050083c8150003c8250083c6350023806700a380170123810701a381d70091059107e30307e283c6050003c715008907238fd7fea38fe7fe890539b513f73700e31d07ec39b59306c6fe93f306ff1384170093841500938213012380170113d94600ae92a687a28803a8370083a5770083a6b7001b53870003a7f7009b1f88011b9f85019b9e86011b5888009bd585009bd686001b1e87013363f3013368e801b3e5d501b3e6c60123a0680023a2080123a4b80023a6d800c107c108e39657fa9307190092073d16b385f40033067640a297a1b593d84800938e18002e88033e88000333080085062334c7012330670041084107e3e5d6ff85089208c695c6973d8a01bb9306c6fe03c8150093f306ff13842700938425009382230123801701a380070113d94600ae92a687a28803a8270083a5670083a6a7001b53070103a7e7009b1f08011b9f05019b9e06011b5808019bd505019bd606011b1e07013363f3013368e801b3e5d501b3e6c60123a0680023a2080123a4b80023a6d800c107c108e39657fa9307190092073916b385f40033067640a29749b3aa8709b919ca0347050083c705007d166317f700050585057df6014582800345050083c705001d9d8280aa862e87b287630db50cb388c5403308c040b388a84006082e832a8e6372181b3346b5001d8a637fb50a63010612cdcb1386f7ff9d4563f8c51813061700b305c54093b5750093c5150093f5f50f638a0516b365e5009d896395051693f587ffba95033603002103210e233ccefee39a65fe13f687ff13f57700aa87b385c600329739cd0345070005462380a5006389c704034517000946a380a5006382c704034527000d462381a500638bc702034537001146a381a5006384c7020345470015462382a500638dc700034557001946a382a5006386c700834767002383f5003685828029ea3306f5001d8a65ca1386f7fffdd7b307c5007d5821a07d16e30106ffb305c70003c5050093f57700fd17a380a700e5f59d4763fac70ab2871d48e117b305f7008861b385f60088e1e369f8fe93777600cdd7fd173306f700834506003386f6002300b600f5b71376750041ca9385f7ffc9d72a867d5821a0fd15e38005f903450700050693777600a30fa6fe0507edf79d4763fcb704938885ff93f888ffa10833051601ba8703b807002106a107233c06ffe31aa6fe469793f77500130617008ddfba9711a005060347f6ff0505a30fe5fee31af6fe36858280cdba3685d5b713061700f9bfb287a5b73285ae8713061700e1f919b73e8625bf2a86be8549bf000000000000cdccccccccccccccd182e6ad7f520e5108c9bcf367e6096a1f6c3e2b8c68059b3ba7ca8485ae67bb6bbd41fbabd9831f2bf894fe72f36e3c79217e1319cde05bf1361d5f3af54fa54b598638d6c56d340101010101010101ff00ff00ff00ff00fffefefefefefefe80808080808080800a0a0a0a0a0a0a0aaf47e17a14ae4701555555555555555533333333333333330f0f0f0f0f0f0f0f01010101010101019a9999999999990100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000a0da0a000000000000100000000000000400000000000000a0ca020000000000001008000000000040000000000000000100000000000000300a010000000000000000000000000030b2020000000000011101250e1305030e10171b0eb44219110155170000023901030e0000032e001101120640186e0e030e3a0b3b053f198701190000042e00110112064018030e3a0b3b05360b3f198701190000052e006e0e030e3a0b3b05200b0000062e001101120640186e0e030e3a0b3b050000072e006e0e030e3a0b3b0b200b0000082e011101120640186e0e030e3a0b3b0b360b0000091d00311311011206580b590b570b00000a1d0031135517580b590b570b00000b1d00311311011206580b5905570b00000c1d0031135517580b5905570b00000d2e006e0e030e3a0b3b0b3f19200b00000e2e011101120640186e0e030e3a0b3b0b3f1900000f1d0131135517580b590b570b0000101d01311311011206580b590b570b0000111d01311311011206580b5905570b0000121d0131135517580b5905570b0000132e006e0e030e3a0b3b053f19200b0000142e011101120640186e0e030e3a0b3b05360b3f190000152e011101120640186e0e030e3a0b3b053f190000162e0111011206401831130000172e0011011206401831130000182e001101120640186e0e030e3a0b3b0b0000192e011101120640186e0e030e3a0b3b0b00001a2e011101120640186e0e030e3a0b3b0500001b2e011101120640186e0e030e3a0b3b05360b3f1987011900001c2e001101120640186e0e030e3a0b3b0b3f1987011900001d2e006e0e030e3a0b3b0b870119200b00001e2e001101120640186e0e030e3a0b3b0b360b3f19870119000000700000000400000000000801752b00001c0060460000000000002b13000000000000000000007011000002742f0000020000000003326e0100000000000e00000001527c4f000064380000010b020002742f000002953f000004406e0100000000000e0000000152190f0000028e010300000000242600000400000000000801752b00001c005a170000880000002b1300000000000000000000a0110000023b1a00000284050000052f0d00009017000002f90501062eb3010000000000020000000152dc350000dd0c000002eb0102ab3f0000029733000005e6380000182500000593030105e6380000182500000593030105e6380000182500000593030105e6380000182500000593030105e63800001825000005930301059a2a00006c2300000593030105eb2c0000d14900000593030105ba3b00006f3a00000593030105770c0000f90300000536050105e638000018250000059303010000025f0d0000029733000005ae420000182500000701040105ae420000182500000701040105ae420000182500000701040105ae420000182500000701040105ae420000182500000701040105b03300008d1800000701040105ff0b0000d537000007010401000005a6000000794a00000273040105fd13000057440000027304010524490000900500000249050105b8080000cc00000002490501050b2a0000f903000002610601000293330000025b130000029034000007fd4b00005429000003d00100027b4100000736140000c8490000038e01078f3e000093330000038901078f3e000093330000038901000002544c0000024f3100000830b3010000000000420100000152fc1600007638000004d3030965000000a0b30100000000000200000004f1360ac61b00000000000004f1150972000000b2b30100000000000200000004f2360ad31b00004000000004f215097f000000fab30100000000000200000004fd360ae01b00007000000004fd1509f300000008b40100000000000200000004fd470b0001000022b4010000000000020000000403011e0b8c00000034b401000000000002000000040701360ced1b0000a0000000040701150b0d01000042b401000000000002000000040701470b1a01000050b401000000000006000000040f0133000002550c000007472d0000c03e000004430107441b0000f204000004430107c1160000b410000004430107aa3000004e2b000004430100022a2b00000d01150000581d000004870100028b4700000dc54a00001d3c0000042a010002761500000efebb010000000000700000000152ef30000093330000049a0fd902000020090000049b11103c1d000004bc01000000000008000000044e1d11a71c000004bc0100000000000800000019f80209094101000004bc010000000000080000001bef5000000a0f0300005009000004511c09ec21000016bc01000000000004000000045116092103000024bc010000000000080000000451280fd824000080090000046514120b1e0000b0090000225901090af81d0000e0090000171209000000000002c60700000d73350000581d000004870100020f0f00000ed6c2010000000000720000000152f528000093330000049a0fe5020000100e0000049b1110901d0000dcc201000000000008000000044e1d11a71c0000dcc20100000000000800000019f802090941010000dcc2010000000000080000001bef5000000afa030000400e000004511c09f9210000f2c20100000000000400000004511609b11b0000fec201000000000008000000044f190fe5240000700e000004651412171e0000a00e0000225901090af81d0000d00e00001712090000000000024b4800000e48c3010000000000720000000152af48000093330000049a0ff1020000000f0000049b11109d1d00004ec301000000000008000000044e1d11a71c00004ec30100000000000800000019f8020909410100004ec3010000000000080000001bef5000000a0f030000300f000004511c090622000064c30100000000000400000004511609b11b000070c301000000000008000000044f190ff2240000600f000004651412231e0000900f0000225901090af81d0000c00f0000171209000000000002210800000e72c40100000000007000000001521f03000093330000049a0ffd02000080100000049b1110aa1d000078c401000000000008000000044e1d11a71c000078c40100000000000800000019f80209094101000078c4010000000000080000001bef5000000afa030000b010000004511c09132200008ac401000000000004000000045116092103000098c4010000000000080000000451280fff240000e0100000046514122f1e000010110000225901090af81d00004011000017120900000000000002d74d000013e90a00001e0b000008bd0601137f0300005331000008f6060113c94c00004344000008100701056b0d000088050000086e05011472b4010000000000e4010000015289020000cc34000008de04030b6206000090b40100000000000c00000008e504130b6f060000acb40100000000000400000008ea04190b7c060000e8b401000000000002000000080a051a1289060000d00000000817052411df1f0000d0b5010000000000040000000880051211cc1f0000d0b5010000000000040000000ec702090b32220000d0b5010000000000020000000e6d020c000000121b13000010010000081a051112ec1f0000400100000894041212cc1f0000700100000ec702090c32220000a00100000e6d020c00000012c8210000d0010000080b05200b5001000062b501000000000006000000139403160b6a01000076b501000000000004000000139503090012d521000000020000080c05210b5d01000068b501000000000004000000139403160b770100007ab5010000000000040000001395030900118906000094b50100000000001a000000080e052411df1f00009ab5010000000000040000000880051211cc1f00009ab5010000000000040000000ec702090b322200009ab5010000000000040000000e6d020c0000001184200000beb40100000000001c00000008eb0416101f200000beb40100000000001c0000001231091013200000beb40100000000001c00000011200910771f0000beb40100000000001c00000011874c10ea1e0000beb40100000000001c000000105331111d1f0000beb40100000000001c0000000a940d09104d1f0000beb40100000000001c0000000c321110dd1e0000beb40100000000001c0000000f7c09120a1c0000300200000ab0091d104c1c0000cab401000000000002000000092b350927010000cab4010000000000020000000953520000125f1f0000800200000ab10915108d1f0000ccb4010000000000080000000f541c1030200000ccb40100000000000800000010501609db200000ccb40100000000000800000011871f0000092e1f0000d6b4010000000000020000000f54150000000000000000000015acb6010000000000780300000152784b0000e5300000083c0512a6220000b0020000083e05170c99220000e00200001483020f001136210000dab601000000000004000000084705251129210000dab6010000000000040000001641033311ba1c0000dab6010000000000040000001608032711581c0000dab60100000000000400000019e502090999000000dab6010000000000040000001b62500000000011041f0000deb6010000000000da0000000847052311f71e0000deb60100000000006e0000000a8b010912a2200000100300000a5801100f9020000040030000128c190fe720000070030000122c12090a1c000002b7010000000000040000000b260e09ff2000001ab7010000000000040000000b3212090b21000026b70100000000000a0000000b391309172100003cb70100000000000a0000000b412509f320000016b7010000000000040000000b2e1000000011f91f0000feb6010000000000040000000a57011211cc1f0000feb6010000000000040000000ec702090b32220000feb6010000000000020000000e6d020c00000011a22000006ab70100000000004e0000000a8c010910902000006ab70100000000004a000000128c1910e72000006ab70100000000004a000000122c12090a1c00006ab7010000000000040000000b260e0917210000a2b70100000000000c0000000b4125090b21000096b7010000000000040000000b391309ff20000092b7010000000000040000000b321200000000124f210000a0030000084c05131274210000d003000016b901091143210000b8b7010000000000120000001814010c10c71c0000beb70100000000000400000016dc1f0bc21d0000beb701000000000004000000195a010f000000000cb322000000040000084c051c1184200000ecb70100000000007201000008590523101f200000ecb7010000000000720100001231091013200000f2b70100000000001e00000011200910771f0000f2b70100000000001e00000011874c10ea1e0000f2b70100000000001e000000105331111d1f0000f2b70100000000001e0000000a940d09104d1f0000f2b70100000000001e0000000c321110dd1e0000f2b70100000000001e0000000f7c09120a1c0000300400000ab0091d104c1c0000feb701000000000002000000092b350927010000feb7010000000000020000000953520000125f1f0000800400000ab10915108d1f000000b8010000000000080000000f541c103020000000b80100000000000800000010501609db20000000b80100000000000800000011871f0000092e1f00000ab8010000000000020000000f541500000000000000103d20000010b80100000000004e01000011220910d41c000010b801000000000014000000113a270b8401000010b80100000000000600000019d60d1f11ee1c000016b80100000000000800000019da0d200be11c000016b80100000000000800000019460617000bfb1c00001eb80100000000000600000019db0d2400101320000024b80100000000001a00000011471510771f000024b80100000000001a00000011874c10ea1e000024b80100000000001a000000105331111d1f000024b80100000000001a0000000a940d09104d1f000024b80100000000001a0000000c321110dd1e000024b80100000000001a0000000f7c09120a1c0000b00400000ab0091d104c1c00002eb801000000000002000000092b3509270100002eb8010000000000020000000953520000125f1f0000000500000ab10915108d1f000030b8010000000000080000000f541c103020000030b80100000000000800000010501609db20000030b80100000000000800000011871f0000092e1f00003ab8010000000000020000000f541500000000000000101320000040b80100000000001c00000011473510771f000040b80100000000001c00000011874c10ea1e000040b80100000000001c000000105331111d1f000040b80100000000001c0000000a940d09104d1f000040b80100000000001c0000000c321110dd1e000040b80100000000001c0000000f7c09120a1c0000300500000ab0091d104c1c00004cb801000000000002000000092b3509270100004cb8010000000000020000000953520000125f1f0000800500000ab10915108d1f00004eb8010000000000080000000f541c10302000004eb80100000000000800000010501609db2000004eb80100000000000800000011871f0000092e1f000058b8010000000000020000000f541500000000000000104920000092b801000000000012000000115a12091f2300009eb801000000000004000000117f0e0010951c0000c0b80100000000000600000011501910151d0000c0b8010000000000060000001b1a0e11641c0000c0b80100000000000600000019e5020909a6000000c0b8010000000000060000001b62500000000a161c0000b00500001150190a55200000f005000011541b0f221c00006006000011631a10701c000032b901000000000002000000092b35093401000032b9010000000000020000000953520000096120000034b90100000000000c00000011641b106d2000004ab901000000000012000000116616092c23000056b901000000000004000000117f0e0009081d0000bcb801000000000004000000114f2c10821c0000a8b801000000000010000000114a121181220000b4b8010000000000040000001bcb051b1173220000b4b8010000000000040000000d7e04080b61220000b4b8010000000000040000000d2e03090000000000001289060000b00600000863052811df1f0000bab9010000000000040000000880051211cc1f0000bab9010000000000040000000ec702090b32220000bab9010000000000020000000e6d020c000000111b130000e6b9010000000000260000000865051512ec1f0000f00600000894041212cc1f0000200700000ec702090c32220000500700000e6d020c000000000d8b3b00000430000008f20113981800003d2d000008f4050113123400001d2b00000843070105c1280000ea1d0000089c04011630c20100000000009800000001520813000011ca1900003cc20100000000001800000008e6071b0b0b1200003cc20100000000000c0000001f17011200116718000062c20100000000005800000008e8070911ac2400006cc20100000000004a0000001f650127115b1700006ec20100000000004800000020270516116f17000082c2010000000000060000001f66013c0b6f06000082c2010000000000060000001f700109000b0b1200008ac2010000000000140000001f6701150b0b120000a0c2010000000000160000001f6901110000000013db070000fe24000008e507010002c51b00000559180000e7310000089304010002ed31000002cc3400000656b6010000000000560000000152874d00007f1b000008f304000005ac090000434d0000086404010517100000d1090000087904011532ba0100000000007e0100000152943c0000e73100000838040cff110000800700000839041912a71f0000b0070000084d041d0a2e1c0000e00700001d2f1100124f130000100800000856041a115c130000baba01000000000018000000086b04150bb3010000c0ba010000000000120000000881042c00115c130000e0ba01000000000018000000086c04190bb3010000e6ba010000000000120000000881042c0011221d000000bb010000000000040000000873041f11ce1d000000bb010000000000040000001996011a09b300000000bb0100000000000400000017ee1c00000bbf01000004bb010000000000080000000876040b0012b31f000040080000083f041d0a3a1c0000700800001d2f11000bcb01000052bb0100000000000a00000008460415122f1d0000a0080000085d042612da1d0000e0080000195a010f10e61d000080bb0100000000000400000017d93609c000000080bb0100000000000400000017ee1c0000000002f101000007244000000c3c00001f5501023b3b00000e6ebc010000000000bc01000001527e3800003d2d00001f1f0fc7200000100a00001f201212b4200000400a0000123f050911b3210000f4bc010000000000d40000001272020f11561d0000febc01000000000008000000249e01320b411e0000febc01000000000008000000195a010900118b1e000006bd010000000000ac00000024a2012209971e00000cbd0100000000001a000000252c1010a31e000026bd0100000000008c000000252f0510cd00000026bd0100000000000c0000002552160b8401000026bd0100000000000c000000054005160010bb1e00006cbd0100000000000a000000256a1609462300006cbd010000000000020000002514070010af1e000056bd0100000000000a000000256916093923000056bd010000000000020000002514070009da0000004abd0100000000000400000025651b09971e00009ebd0100000000001400000025771609971e00007ebd01000000000012000000255a1e000011631d0000bebd0100000000000200000024b701430b411e0000bebd01000000000002000000195a0109001152220000c0bd0100000000000400000024b8011c11781e0000c0bd010000000000040000000da9050d095a1e0000c0bd01000000000004000000231a0900000000000f5c210000700a00001f252712a0210000a00a0000165f040d128d210000d00a00002445022912491d0000000b000024de03091145220000d0bc0100000000000a00000019090913116c1e0000d0bc0100000000000a0000000da9050d095a1e0000d0bc0100000000000a000000231a09000000000000000002b140000002454800000592040000542900001f35010100023d1b000005a3240000542900001f650101000002432b000005474d0000664a00001f6f01011510c00100000000002001000001526f0a0000454800001f34011292240000b00b00001f350123114817000034c0010000000000de00000020270516126f170000e00b00001f3601100c6f060000100c00001f700109000b0b1200005cc0010000000000160000001f3801150c0b120000400c00001f4101110bbf24000092c0010000000000020000001f410111127a180000700c00001f3c01220f25120000b00c00001f1a091191180000b2c00100000000000a00000008a3041209c0220000b2c00100000000000a0000001f1a260000000b0b120000fec0010000000000120000001f3e011100000013641e00003d1b00001f63010100026d4b000007291e00000f3000001f15010002a3090000020f300000070b380000542900001f1a01000002321b00000514300000ec0400001f7b010105cf0e0000664a00001f9101010002114d000002ec0400000550300000542900001f7c0101000002dc3a00001530c10100000000000001000001524b050000ec0400001fd40112a4180000f00c00001fd50109129f240000200d00001f7c012311c91800006cc1010000000000c40000002027051612b1180000500d00001f7d01100c6f060000800d00001f920109000b0b12000080c1010000000000180000001f8801150b0b120000a6c1010000000000180000001f7f0115127a180000b00d00001f8301220f25120000e00d00001f1a091191180000d2c10100000000000a00000008a3041209c0220000d2c10100000000000a0000001f1a260000000b0b1200001ac2010000000000160000001f85011100000000000555340000932400001f1301010002d4320000162abe010000000000b400000001523c1a0000101626000038be0100000000009600000008a41a110426000038be010000000000960000002679022a0cf7250000300b000026b6060f00000017debe010000000000380000000152481a000007ae190000da32000008a3010714480000514f000008bf010002973300001816bf0100000000000a0000000152a74b00007745000008c61920bf010000000000b60000000152a2450000da32000008ca103c1a00002ebf010000000000a200000008cb09101626000030bf0100000000009600000008a41a110426000030bf010000000000960000002679022a0cf7250000700b000026b6060f0000000019d6bf0100000000003a0000000152e53a0000514f000008ce09481a0000f6bf0100000000001400000008cf090000022a0a000005da1000009333000008bb09010002d30c00001abac30100000000001600000001524b3300002511000008d0080b0e1b0000bac30100000000001600000008d0083e00000002db3c000002ce4d0000024d4c0000192ab3010000000000040000000152340a0000b54f000001fa10a10100002ab30100000000000400000001fa0509340000002ab30100000000000200000003d21e0000000002242f000002d0070000052a2f0000b01000002742020100000002df3c000005ab0a00008e110000065f0a0105ab0a00008e110000065f0a0105ab0a00008e110000065f0a0105ab0a00008e110000065f0a0100029d34000002a11e0000022025000007663600000e490000097c0107153e0000c1010000097c0107712c000076440000097c01076b4e00005a410000097c0107a01c000006400000097c010002383900000712000000a41b0000094b0107812f0000094d00001b5b0107e13400007c2300001b5b01078c2300004b370000094b010002614e000005ef390000764400001bc7050100029733000007740b0000ff3d00001b190100024d0c0000071a1d00002c4500001bd90100000297330000058a120000d11b000019e4020105501c0000fc2900001956010105404700009a4a000019cb0d01052c270000fb400000199806010518060000124100001942060105924400006209000019860d01053a2a0000862a00001916040105443b0000ee3d000019e4020105b41a0000d1120000198f010105e64400002f3200001956010105c6270000da09000019f70201055b0e00002b19000019040901054c0400000a1b000019560101054c0400000a1b00001956010102b607000003c8c20100000000000e0000000152fa450000c93c0000190b0d0005c6270000da09000019f7020105c6270000da09000019f7020105c6270000da09000019f702010002b4030000023b3b000007af050000d934000017d7010761370000f62a000017e30107f20d0000ff12000017d7010784410000fe33000017e3010002793a000005fa010000ee49000017ec01010002973300000740320000cd1800001711010740320000cd1800001711010740320000cd1800001711010740320000cd1800001711010002b140000005e9150000d9340000175f01010000029e0d000002114d00000780150000e73e0000235201000297330000075e1d0000a6400000231901075e1d0000a64000002319010000020830000007391900000830000025290107f53e00002d3f00002534010d2c4b0000db1d00002547010772100000f84100002513010772100000f8410000251301000002a11e0000027a2f000002b62b00000298460000055e1300002b2500000aaa090105b53f0000fc4200000a8f0d01057b390000f60000000a56010105ec080000b60f00000a8a0101000002a611000002ac1100000760290000ea3c00000c310102670d000007cf430000b61100000c35010000000002704a0000025d310000023b3b00000761310000a61e00000f78010002e84d000007ad460000c32000000f5401000002e14d0000023b3b0000072b0800009e130000104d01020c000000021749000007a5170000590000001050010000000002961c000002a30900000763060000822700001d2e01076c140000d32300001d2e0100000002df080000023b3b0000054b490000712200000e6c02010002844a00000582220000764400000ec602010582220000764400000ec602010582220000764400000ec602010000000208000000020c0000000d280b00008c1b000011860107230f0000a1460000111a01028c1b0000076520000054290000118701000d2b090000a51a0000112601071f41000023140000117a01072a2c0000d2010000117201072a2c0000d2010000117201071f41000023140000117a010002a11e0000029733000007584c00000c00000012300107f14d00001f0100001229010002114d000007da1b00001f010000128a010002bb3200000517280000620c0000126c020100025a45000005e82d0000c9320000123e0501000002680b000007ba400000f43f00000b180107bf2b0000c23900000b240107d80f0000fe2b00000b0b010717230000592300000b11010717230000592300000b11010717230000592300000b1101000297330000053d390000e33600001607030105b62900008d4a00001640030107a80d00000e2c000016d30105e93600002537000016b80101050a04000096400000165b040100027a2f000002a73300000524010000ab05000018130101000002174b0000022a2b000005e54e00001f4b000024dd03010002844a000005652800001f4b000024410201000297330000056a2e000026350000249b0101000000022049000005b63d0000b71b0000138f030105a3340000570f0000138f030102822d0000026a15000005bd470000bb4a000021e8010105bd470000bb4a000021e8010105bd470000bb4a000021e8010105bd470000bb4a000021e80101000000029e0d000002a20d000002ec00000005401a0000e03600000d53050100028a24000005233c0000342b00000da8050105233c0000342b00000da8050100000595470000f63100000d930401026b3a0000051a4d00001f2c00000d2a030100057e0900001f2c00000d7d04010002e508000002a033000005790f00009c050000145602010503470000df3d00001482020105ba0300008244000014bb030105f6060000a70e000014120601001be2bb0100000000000e00000001527b420000bb3c0000148b0703117f230000e4bb0100000000000c000000148c07050973230000e4bb0100000000000c0000001c860500000002544c0000028b47000005bc2f0000ae4a00001ae4040105bc2f0000ae4a00001ae40401051e4a0000444f00001acd0401051e4a0000444f00001acd0401000002ec2a00001c24ba0100000000000e00000001522d170000e93000001c6e1d60400000091300001c95011d411000004b3400001c85011ef0bb0100000000000e000000015210330000644500001c50030002051b000002bc27000015b0bb01000000000012000000015255480000933300001ebb021118120000b0bb010000000000120000001ebc021b11dd140000b0bb0100000000001200000008440709090b120000b0bb010000000000120000001f591200000000021c35000015c2bb010000000000120000000152c2020000933300001ed6021118120000c2bb010000000000120000001ed7021b11dd140000c2bb0100000000001200000008440709090b120000c2bb010000000000120000001f5912000000000002fa14000003d4bb0100000000000e0000000152180500001d13000020720602664b00000531350000e1190000202505010532070000823a00002025050105740700003a3f000020250501000206330000050b4200000d0a0000209b0701000002112800000221190000050a2400008f2d000022580101050a2400008f2d000022580101050a2400008f2d000022580101050a2400008f2d0000225801010002063300000ed0c3010000000000a200000001522d1100009333000022830f08130000f00f000022830a12ca1900002010000008e6071b0c0b120000501000001f1701120011671800000ec40100000000005800000008e8070911ac24000018c40100000000004a0000001f650127115b1700001ac40100000000004800000020270516116f1700002ec4010000000000060000001f66013c0b6f0600002ec4010000000000060000001f700109000b0b12000036c4010000000000140000001f6701150b0b1200004cc4010000000000160000001f6901110000000000000002f1060000020338000005e12e00006a190000269906010573190000142f000026b5060102973300000572160000084800002677020100000000003c0000000200000000000800ffffffff326e0100000000000e00000000000000406e0100000000000e0000000000000000000000000000000000000000000000ec0100000200740000000800ffffffff2ab301000000000004000000000000002eb3010000000000020000000000000030b3010000000000420100000000000072b4010000000000e40100000000000056b60100000000005600000000000000acb6010000000000780300000000000024ba0100000000000e0000000000000032ba0100000000007e01000000000000b0bb0100000000001200000000000000c2bb0100000000001200000000000000d4bb0100000000000e00000000000000e2bb0100000000000e00000000000000f0bb0100000000000e00000000000000febb01000000000070000000000000006ebc010000000000bc010000000000002abe010000000000b400000000000000debe010000000000380000000000000016bf0100000000000a0000000000000020bf010000000000b600000000000000d6bf0100000000003a0000000000000010c0010000000000200100000000000030c1010000000000000100000000000030c20100000000009800000000000000c8c20100000000000e00000000000000d6c2010000000000720000000000000048c30100000000007200000000000000bac30100000000001600000000000000d0c3010000000000a20000000000000072c4010000000000700000000000000000000000000000000000000000000000a2b3010000000000a6b3010000000000aab3010000000000b2b3010000000000beb3010000000000c2b301000000000000000000000000000000000000000000b4b3010000000000bcb3010000000000c2b3010000000000cab301000000000000000000000000000000000000000000fcb301000000000008b40100000000000ab401000000000014b40100000000000000000000000000000000000000000036b401000000000042b401000000000044b40100000000004cb401000000000000000000000000000000000000000000ecb4010000000000f2b4010000000000f6b4010000000000fcb4010000000000b0b5010000000000e0b50100000000000000000000000000000000000000000010b601000000000030b601000000000050b601000000000056b60100000000000000000000000000000000000000000018b601000000000020b601000000000050b601000000000056b60100000000000000000000000000000000000000000018b601000000000020b601000000000050b601000000000056b60100000000000000000000000000000000000000000018b601000000000020b601000000000050b601000000000056b60100000000000000000000000000000000000000000062b501000000000068b501000000000076b50100000000007ab50100000000000000000000000000000000000000000068b50100000000006cb50100000000007ab50100000000007eb501000000000000000000000000000000000000000000beb4010000000000c2b4010000000000cab4010000000000ccb4010000000000d4b4010000000000d6b4010000000000d8b4010000000000dab401000000000000000000000000000000000000000000ccb4010000000000d4b4010000000000d6b4010000000000d8b401000000000000000000000000000000000000000000aeb6010000000000c4b6010000000000c6b6010000000000ceb601000000000000000000000000000000000000000000aeb6010000000000c4b6010000000000c6b6010000000000ceb601000000000000000000000000000000000000000000f0b6010000000000fab601000000000002b70100000000004cb701000000000000000000000000000000000000000000f0b6010000000000f4b601000000000002b701000000000048b701000000000000000000000000000000000000000000f0b6010000000000f4b601000000000002b701000000000048b701000000000000000000000000000000000000000000b8b7010000000000ceb7010000000000d4b7010000000000d8b701000000000000000000000000000000000000000000b8b7010000000000ceb7010000000000d4b7010000000000d8b701000000000000000000000000000000000000000000d0b7010000000000d4b7010000000000dab7010000000000dcb701000000000000000000000000000000000000000000f2b7010000000000f6b7010000000000feb701000000000000b801000000000008b80100000000000ab80100000000000cb801000000000010b80100000000000000000000000000000000000000000000b801000000000008b80100000000000ab80100000000000cb80100000000000000000000000000000000000000000024b801000000000028b80100000000002eb801000000000030b801000000000038b80100000000003ab80100000000003cb80100000000003eb80100000000000000000000000000000000000000000030b801000000000038b80100000000003ab80100000000003cb80100000000000000000000000000000000000000000040b801000000000042b80100000000004cb80100000000004eb801000000000056b801000000000058b80100000000005ab80100000000005cb8010000000000000000000000000000000000000000004eb801000000000056b801000000000058b80100000000005ab801000000000000000000000000000000000000000000c6b8010000000000c8b80100000000000cb901000000000010b901000000000012b901000000000018b901000000000000000000000000000000000000000000d0b8010000000000d8b8010000000000dab8010000000000deb8010000000000e0b8010000000000e6b8010000000000e8b8010000000000f8b8010000000000fab8010000000000fcb801000000000000b90100000000000cb90100000000000000000000000000000000000000000018b901000000000030b901000000000032b901000000000034b901000000000040b901000000000042b901000000000044b901000000000048b90100000000000000000000000000000000000000000062b901000000000068b90100000000006cb901000000000072b901000000000098b9010000000000cab901000000000000000000000000000000000000000000eeb9010000000000f6b901000000000008ba0100000000000cba01000000000000000000000000000000000000000000eeb9010000000000f6b901000000000008ba0100000000000cba01000000000000000000000000000000000000000000eeb9010000000000f2b901000000000008ba0100000000000cba010000000000000000000000000000000000000000004aba01000000000052ba01000000000056ba0100000000005eba0100000000000000000000000000000000000000000064ba0100000000008eba0100000000000ebb0100000000001ebb0100000000000000000000000000000000000000000064ba0100000000008eba0100000000000ebb0100000000001ebb01000000000000000000000000000000000000000000a0ba010000000000aeba010000000000b2ba0100000000000cbb0100000000000000000000000000000000000000000022bb01000000000040bb0100000000005ebb01000000000068bb0100000000000000000000000000000000000000000022bb01000000000040bb0100000000005ebb01000000000068bb010000000000000000000000000000000000000000006cbb01000000000072bb01000000000078bb0100000000007cbb01000000000080bb01000000000084bb010000000000000000000000000000000000000000006cbb01000000000072bb01000000000078bb0100000000007cbb01000000000080bb01000000000084bb0100000000000000000000000000000000000000000004bc0100000000005abc01000000000060bc0100000000006ebc0100000000000000000000000000000000000000000014bc01000000000016bc0100000000002cbc01000000000030bc010000000000000000000000000000000000000000003abc01000000000044bc01000000000060bc0100000000006ebc010000000000000000000000000000000000000000003abc01000000000044bc01000000000060bc0100000000006ebc010000000000000000000000000000000000000000003abc01000000000044bc01000000000060bc0100000000006ebc01000000000000000000000000000000000000000000b4bc010000000000ccbc010000000000ecbc010000000000c8bd01000000000000000000000000000000000000000000b4bc010000000000ccbc010000000000ecbc010000000000c8bd01000000000000000000000000000000000000000000ccbc010000000000dabc010000000000f8bd010000000000fcbd01000000000000000000000000000000000000000000ccbc010000000000dabc010000000000f8bd010000000000fcbd01000000000000000000000000000000000000000000ccbc010000000000dabc010000000000f8bd010000000000fcbd01000000000000000000000000000000000000000000ccbc010000000000dabc010000000000f8bd010000000000fcbd0100000000000000000000000000000000000000000038be0100000000003cbe01000000000044be0100000000004abe01000000000066be0100000000006cbe0100000000000000000000000000000000000000000030bf01000000000034bf0100000000003cbf01000000000042bf0100000000005ebf01000000000064bf0100000000000000000000000000000000000000000026c001000000000028c001000000000034c001000000000012c10100000000000000000000000000000000000000000038c00100000000003cc001000000000040c001000000000044c00100000000000000000000000000000000000000000038c00100000000003cc001000000000040c001000000000044c00100000000000000000000000000000000000000000082c00100000000008cc00100000000008ec001000000000092c001000000000000000000000000000000000000000000a0c0010000000000a4c0010000000000aac0010000000000e8c0010000000000ecc0010000000000f6c001000000000000000000000000000000000000000000a0c0010000000000a4c0010000000000aac0010000000000e8c0010000000000ecc0010000000000f6c00100000000000000000000000000000000000000000042c101000000000054c10100000000006cc101000000000030c2010000000000000000000000000000000000000000004ac10100000000004cc10100000000006cc101000000000030c20100000000000000000000000000000000000000000070c101000000000074c101000000000078c10100000000007cc10100000000000000000000000000000000000000000070c101000000000074c101000000000078c10100000000007cc101000000000000000000000000000000000000000000c0c1010000000000c4c1010000000000cac101000000000012c201000000000000000000000000000000000000000000c0c1010000000000c4c1010000000000cac101000000000012c201000000000000000000000000000000000000000000dcc201000000000034c30100000000003ac301000000000048c301000000000000000000000000000000000000000000f0c2010000000000f2c201000000000006c30100000000000ac30100000000000000000000000000000000000000000014c30100000000001ec30100000000003ac301000000000048c30100000000000000000000000000000000000000000014c30100000000001ec30100000000003ac301000000000048c30100000000000000000000000000000000000000000014c30100000000001ec30100000000003ac301000000000048c3010000000000000000000000000000000000000000004ec3010000000000a6c3010000000000acc3010000000000bac30100000000000000000000000000000000000000000062c301000000000064c301000000000078c30100000000007cc30100000000000000000000000000000000000000000086c301000000000090c3010000000000acc3010000000000bac30100000000000000000000000000000000000000000086c301000000000090c3010000000000acc3010000000000bac30100000000000000000000000000000000000000000086c301000000000090c3010000000000acc3010000000000bac301000000000000000000000000000000000000000000dac3010000000000dcc3010000000000dec301000000000066c401000000000000000000000000000000000000000000dac3010000000000dcc3010000000000dec3010000000000fac301000000000000000000000000000000000000000000dac3010000000000dcc3010000000000dec3010000000000eec30100000000000000000000000000000000000000000078c4010000000000cec4010000000000d4c4010000000000e2c40100000000000000000000000000000000000000000088c40100000000008ac4010000000000a0c4010000000000a4c401000000000000000000000000000000000000000000aec4010000000000b8c4010000000000d4c4010000000000e2c401000000000000000000000000000000000000000000aec4010000000000b8c4010000000000d4c4010000000000e2c401000000000000000000000000000000000000000000aec4010000000000b8c4010000000000d4c4010000000000e2c401000000000000000000000000000000000000000000326e010000000000406e010000000000406e0100000000004e6e010000000000000000000000000000000000000000002ab30100000000002eb30100000000002eb301000000000030b301000000000030b301000000000072b401000000000072b401000000000056b601000000000056b6010000000000acb6010000000000acb601000000000024ba01000000000024ba01000000000032ba01000000000032ba010000000000b0bb010000000000b0bb010000000000c2bb010000000000c2bb010000000000d4bb010000000000d4bb010000000000e2bb010000000000e2bb010000000000f0bb010000000000f0bb010000000000febb010000000000febb0100000000006ebc0100000000006ebc0100000000002abe0100000000002abe010000000000debe010000000000debe01000000000016bf01000000000016bf01000000000020bf01000000000020bf010000000000d6bf010000000000d6bf01000000000010c001000000000010c001000000000030c101000000000030c101000000000030c201000000000030c2010000000000c8c2010000000000c8c2010000000000d6c2010000000000d6c201000000000048c301000000000048c3010000000000bac3010000000000bac3010000000000d0c3010000000000d0c301000000000072c401000000000072c4010000000000e2c4010000000000000000000000000000000000000000007261775f7665630073747200636f756e74005f5a4e34636f726535736c6963653469746572313349746572244c542454244754243134706f73745f696e635f73746172743137683231633736663939343638653065646545007b636c6f7375726523307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e005f5a4e34636f726533707472347265616431376831626239643039646638396234373532450077726974653c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e007b696d706c2335347d00616476616e63655f62793c636f72653a3a7374723a3a697465723a3a43686172496e64696365733e006e657874005f5a4e34636f726533737472367472616974733131305f244c5424696d706c2475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c5424737472244754242475323024666f722475323024636f72652e2e6f70732e2e72616e67652e2e52616e6765546f244c54247573697a652447542424475424336765743137683633326532303137643665353735396645006e6578743c5b7573697a653b20345d3e00636f6e7461696e735f6e6f6e5f636f6e74696e756174696f6e5f62797465006275696c64657273005f5a4e3131305f244c5424636f72652e2e6f70732e2e72616e67652e2e52616e676546726f6d244c54247573697a6524475424247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c54242475356224542475356424244754242447542435696e6465783137686163396536316662616530626263376145005f5a4e34636f726533666d7439466f726d617474657231327061645f696e74656772616c3137686238656639343965396131613633346545005f5a4e36335f244c5424636f72652e2e63656c6c2e2e426f72726f774d75744572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683636336332373865383138373636393045005f5a4e34636f726533666d74336e756d35335f244c5424696d706c2475323024636f72652e2e666d742e2e55707065724865782475323024666f7224753230246936342447542433666d743137683464336136353331313038303933376445005f5a4e34636f726533666d7439466f726d617474657239616c7465726e617465313768333537326537646636323036356664374500696e646578005f5a4e34636f7265366f7074696f6e31354f7074696f6e244c5424542447542439756e777261705f6f72313768343165333439646137383638346138334500616c69676e5f6f66667365743c75383e005f5a4e34636f72653373747232315f244c5424696d706c24753230247374722447542439656e64735f776974683137683139626662313333653233336465306145005f5a4e34636f726535736c69636532395f244c5424696d706c2475323024247535622454247535642424475424336765743137683233646638653962656438656665346645005f5a4e34636f726533666d74386275696c64657273313044656275675475706c65356669656c6432385f24753762242475376224636c6f7375726524753764242475376424313768636364396362623165623562613563364500656e74727900666d745f696e743c636f72653a3a666d743a3a6e756d3a3a55707065724865782c2075383e005f5a4e34636f726536726573756c743133756e777261705f6661696c65643137683030653934303161326339653536633045005f5a4e34636f726533666d74386275696c6465727338446562756753657435656e7472793137686531623638303262326163636539656445007074720070616464696e670077726974653c636861723e0069735f736f6d653c7573697a653e00676574005f5a4e37355f244c54247573697a65247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c542424753562245424753564242447542424475424336765743137683362336666656535366439303731313345005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243873706c69745f61743137683461343239666364306233623563343945005f5a4e3131305f244c5424636f72652e2e697465722e2e61646170746572732e2e656e756d65726174652e2e456e756d6572617465244c54244924475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e65787431376831623734616564656639323065303665450063686172005f5a4e34636f7265366f7074696f6e31354f7074696f6e244c5424542447542436696e736572743137686265366237313331636461646331646245005f5a4e34636f726536726573756c743139526573756c74244c542454244324452447542438616e645f7468656e3137683138643933303364393238646565393245005f5a4e34636f726536726573756c743139526573756c74244c542454244324452447542438616e645f7468656e313768316532623263316238653933626561654500636f70795f66726f6d5f736c696365007b696d706c2332397d007b696d706c233232357d005f5a4e34636f726533666d7439466f726d6174746572323564656275675f7475706c655f6669656c64315f66696e6973683137683963326264643732306464613133376545007b696d706c2336357d005f5a4e3130385f244c5424636f72652e2e697465722e2e61646170746572732e2e66696c7465722e2e46696c746572244c5424492443245024475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722447542435636f756e743137683631323362313132363938303130326445005f5a4e34636f72653370747235777269746531376830336462313664353065636536366165450072616e6765006f7074696f6e005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f72336e74683137683635613666633036633265613031396645005f5a4e34636f72653373747235636f756e743134646f5f636f756e745f6368617273313768653066306166323562653730356463664500616c69676e5f746f5f6f6666736574733c75382c207573697a653e005f5a4e34636f726533636d70336d696e3137683961303232643031326665326338333745007b696d706c23317d005f5a4e34636f726533666d743372756e313768666639613633333362396633663061614500676574636f756e7400697465725f6d75743c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e006272616e63683c28292c20636f72653a3a666d743a3a4572726f723e007b696d706c2332357d005f5a4e34636f7265336f70733866756e6374696f6e36466e4f6e63653963616c6c5f6f6e63653137683331326365396462383432326365623645005f5a4e34636f726533666d74386275696c64657273313044656275675475706c65356669656c643137686134393061356537663734366534656245005f5a4e34636f72653130696e7472696e736963733139636f70795f6e6f6e6f7665726c617070696e673137683165326664363834393232323263326345005f5a4e34636f726533666d7439466f726d6174746572397369676e5f706c75733137683765363563323535316433616561343445007369676e5f706c7573005f5a4e34636f72653373747235636f756e743233636861725f636f756e745f67656e6572616c5f6361736531376864313333363866323830386530613030450076616c69646174696f6e73005f5a4e34636f726535736c696365346974657238375f244c5424696d706c2475323024636f72652e2e697465722e2e7472616974732e2e636f6c6c6563742e2e496e746f4974657261746f722475323024666f7224753230242452462424753562245424753564242447542439696e746f5f697465723137683765326332623733366531386264656545005f5a4e34636f726533707472376d75745f70747233315f244c5424696d706c2475323024244250246d75742475323024542447542433616464313768333939313037663564323335643062374500497465724d75740047656e657269635261646978006e6578745f696e636c75736976653c636861723e005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243132616c69676e5f6f66667365743137686265366661383332613635626436303545007b696d706c2335337d0064726f705f696e5f706c6163653c26636f72653a3a697465723a3a61646170746572733a3a636f706965643a3a436f706965643c636f72653a3a736c6963653a3a697465723a3a497465723c75383e3e3e005f5a4e34636f7265337074723133726561645f766f6c6174696c653137683034656338646164326362346562306245006d75745f7074720073756d005f5a4e34636f726533666d7439466f726d61747465723770616464696e67313768386664646163386139653836623737364500636d7000696d706c73005f5a4e34636f72653373747232315f244c5424696d706c247532302473747224475424313669735f636861725f626f756e646172793137683034353265303532643135616334353245005f5a4e37355f244c54247573697a65247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c542424753562245424753564242447542424475424336765743137686337356165633633323166633531643545005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542439656e64735f77697468313768383363653331633938643238356662364500696e736572743c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e005f5a4e34636f726533666d74386275696c6465727331304465627567496e6e65723969735f7072657474793137683430666266303734623763353466303545007b696d706c2334317d005f5f72646c5f6f6f6d005f5a4e34636f72653373747235636f756e743131636f756e745f63686172733137683362393037393633646461313835376345007265706c6163653c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e005f5a4e34636f7265366f7074696f6e31354f7074696f6e244c542454244754243769735f736f6d653137686166353061376333383437653666373645006e74683c636f72653a3a7374723a3a697465723a3a43686172496e64696365733e005f5a4e34636f726533737472313176616c69646174696f6e733135757466385f66697273745f627974653137683962396637633933306431356335663945005f5a4e34636f726533666d7438676574636f756e743137683639663830313763343363306364653245005f5a4e34636f72653970616e69636b696e673970616e69635f7374723137683666303932373830653338346562353045005f5a4e34636f726535736c696365366d656d6368723138636f6e7461696e735f7a65726f5f6279746531376861303536386565313833303061353732450072656d00666d745f696e743c636f72653a3a666d743a3a6e756d3a3a4c6f7765724865782c2075383e005f5a4e34355f244c5424244c502424525024247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d74313768613430323766643039663261636331324500666d743c28293e005f5a4e36375f244c5424636f72652e2e61727261792e2e54727946726f6d536c6963654572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d74313768353264643636336235383463633535664500636f70795f6e6f6e6f7665726c617070696e673c75383e00616363756d007b696d706c2334387d007b636c6f7375726523307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542434697465723137686266616536663139613561623764656445006765745f756e636865636b65643c636f72653a3a666d743a3a72743a3a417267756d656e742c207573697a653e006765743c267374723e0070616e69635f646973706c61793c267374723e00756e777261705f6661696c6564002f72757374632f32663662633564323539653761623235646466646433336465353362383932373730323138393138007274005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f7234666f6c64313768623061333862663336373733633236364500636f756e743c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e005f5a4e34636f726533707472347265616431376831653634383335653639376533366630450073756d5f62797465735f696e5f7573697a65005f5a4e34636f726533666d7432727438417267756d656e743861735f7573697a653137686437613231613332353662616362386245005f5a4e3131305f244c5424636f72652e2e697465722e2e61646170746572732e2e656e756d65726174652e2e456e756d6572617465244c54244924475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e657874313768633030313137313163643937383139624500726573756c74005f5a4e37335f244c5424636f72652e2e666d742e2e6e756d2e2e4c6f776572486578247532302461732475323024636f72652e2e666d742e2e6e756d2e2e47656e657269635261646978244754243564696769743137686634306237613733623764393162653445004d61796265556e696e6974007b696d706c2336347d005f5a4e37335f244c54242475356224412475356424247532302461732475323024636f72652e2e736c6963652e2e636d702e2e536c6963655061727469616c4571244c542442244754242447542435657175616c3137686637383434376536346661643333376145005f5a4e3130365f244c5424636f72652e2e6f70732e2e72616e67652e2e52616e6765244c54247573697a6524475424247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c542424753562245424753564242447542424475424336765743137683761383664333261616263343034303345005f5a4e34636f72653463686172376d6574686f647332325f244c5424696d706c247532302463686172244754243131656e636f64655f757466383137683661333732316366346263313738623645005f5a4e34636f726533666d74336e756d313247656e65726963526164697837666d745f696e743137686363663535643038613665313532386645005f5a4e34636f726533666d74336e756d33696d7037666d745f7536343137683238366534643532373433386334363745005f5a4e34636f72653970616e69636b696e673570616e69633137686437373538656430613265383739363145006c6962726172792f636f72652f7372632f6c69622e72732f402f636f72652e353431663036343835316338633866372d6367752e3000726561645f766f6c6174696c653c7573697a653e005f5a4e3130385f244c5424636f72652e2e697465722e2e61646170746572732e2e66696c7465722e2e46696c746572244c5424492443245024475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722447542435636f756e7438746f5f7573697a6532385f24753762242475376224636c6f73757265247537642424753764243137686532646263323632336436376436643345005f5a4e34636f726533666d743131506f737450616464696e673577726974653137683130373832303864313037663934393045006164643c7573697a653e005f5a4e34636f726533666d7439466f726d61747465723977726974655f737472313768353330393765363135313339346565644500696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e2c20636f72653a3a6f70733a3a72616e67653a3a52616e676546726f6d3c7573697a653e3e007b696d706c2331357d00656e64735f776974683c75383e005f5a4e34636f726535736c696365366d656d636872366d656d6368723137683838333063653264646237323666636245006c656e5f75746638005f5a4e34636f72653463686172376d6574686f64733135656e636f64655f757466385f7261773137686230336466376165346464366562316445005f5a4e34636f726533666d74355772697465313077726974655f63686172313768666466623438666364333637346132384500616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23347d3a3a6669656c643a3a7b636c6f737572655f656e7623307d3e00636f7265005f5a4e34636f726533636d7035696d706c7335375f244c5424696d706c2475323024636f72652e2e636d702e2e5061727469616c4f72642475323024666f7224753230247573697a6524475424326c74313768383563303932356636663163316566654500646f5f636f756e745f6368617273005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542431336765745f756e636865636b656431376838333832313033623533356331333034450063656c6c006765743c75382c20636f72653a3a6f70733a3a72616e67653a3a52616e67653c7573697a653e3e004465627567496e6e65720066696e697368005f5a4e34636f726533666d74336e756d313247656e65726963526164697837666d745f696e7431376835383366363662653034373931303631450077726974655f70726566697800636861725f636f756e745f67656e6572616c5f6361736500706f73745f696e635f73746172743c75383e007265706c6163653c636861723e00506f737450616464696e6700697465723c75383e005f5a4e38375f244c5424636f72652e2e7374722e2e697465722e2e43686172496e6469636573247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683862646365633661316137393933386345005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542433676574313768396431656137353833353464396166364500656e756d6572617465005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683563636236663439653430616432356245005f5a4e34636f726535736c69636534697465723136497465724d7574244c54245424475424336e65773137683131393134666634646337396132326545006469676974005f5a4e34636f726535736c69636533636d7038315f244c5424696d706c2475323024636f72652e2e636d702e2e5061727469616c4571244c54242475356224422475356424244754242475323024666f7224753230242475356224412475356424244754243265713137683331383339323064643563373930336445006d656d6368725f616c69676e656400777261705f6275663c636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23317d3a3a777261703a3a7b636c6f737572655f656e7623307d3e005f5a4e34636f726533666d74386275696c6465727331305061644164617074657234777261703137686630613261643433323636313138356545005f5a4e34636f726533666d74386275696c64657273313044656275675475706c653666696e6973683137683262326465366164386361323965353845006974657200666f6c643c7573697a652c20636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c207573697a652c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e005f5a4e34636f72653373747235636f756e743233636861725f636f756e745f67656e6572616c5f6361736532385f24753762242475376224636c6f73757265247537642424753764243137686238333838383631636166343538396545007b636c6f7375726523307d3c2675382c207573697a652c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e00737065635f6e6578743c7573697a653e005f5a4e34636f726534697465723572616e67653130315f244c5424696d706c2475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722475323024666f722475323024636f72652e2e6f70732e2e72616e67652e2e52616e6765244c5424412447542424475424346e6578743137683166316635393732633862353338396245005f5a4e34636f726533737472313176616c69646174696f6e733138757466385f6163635f636f6e745f62797465313768386431353839303565613233346333334500757466385f6163635f636f6e745f62797465006164643c5b7573697a653b20345d3e006e65773c5b7573697a653b20345d3e005f5a4e34636f726535736c6963653469746572313349746572244c542454244754243134706f73745f696e635f73746172743137686632323465323937613136633263656145006e6578743c636f72653a3a736c6963653a3a697465723a3a497465723c636f72653a3a666d743a3a72743a3a417267756d656e743e3e005f5a4e34636f726535617272617938355f244c5424696d706c2475323024636f72652e2e6f70732e2e696e6465782e2e496e646578244c542449244754242475323024666f722475323024247535622454247533622424753230244e24753564242447542435696e6465783137683663646534633833393961376530333445007b696d706c23397d0064656275675f7475706c655f6e6577005f5a4e34636f726533666d74386275696c64657273313044656275675475706c653666696e69736832385f24753762242475376224636c6f737572652475376424247537642431376861393666623161373161643166373535450064656275675f7475706c655f6669656c64315f66696e697368006164643c75383e007b696d706c233138317d00666f6c643c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a6d61703a3a6d61705f666f6c643a3a7b636c6f737572655f656e7623307d3c2675382c207573697a652c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e3e005f5a4e34636f726535736c69636532395f244c5424696d706c2475323024247535622454247535642424475424313873706c69745f61745f756e636865636b65643137683765396534313435376636393734393145006e6578743c636f72653a3a736c6963653a3a697465723a3a497465723c636f72653a3a666d743a3a72743a3a506c616365686f6c6465723e3e007b696d706c2331377d005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542438697465725f6d75743137683030376635633136366631613761373245006172726179005f5a4e34636f7265337374723469746572323253706c6974496e7465726e616c244c5424502447542431346e6578745f696e636c75736976653137683938613230353930343932666138366445005f5a4e35325f244c542463686172247532302461732475323024636f72652e2e7374722e2e7061747465726e2e2e5061747465726e24475424313269735f7375666669785f6f663137683866653837336364343736333664316445005f5a4e34636f726533666d7439466f726d617474657238777261705f6275663137686636336162363038633262616362303045005f5a4e34636f726533666d74336e756d35325f244c5424696d706c2475323024636f72652e2e666d742e2e55707065724865782475323024666f72247532302469382447542433666d743137683438643832613435336137306166353745007b636c6f7375726523307d005f5a4e35365f244c54247573697a65247532302461732475323024636f72652e2e697465722e2e7472616974732e2e616363756d2e2e53756d244754243373756d3137683739356164323965353439386433333445005f5a4e34636f72653373747232315f244c5424696d706c2475323024737472244754243132636861725f696e64696365733137686466343535663065643137623532303045006765743c75382c207573697a653e005f5a4e34636f7265337074723132616c69676e5f6f66667365743137683534623332333739346162326331313545005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243961735f6368756e6b7331376831643562356538303063366463326238450061735f6368756e6b733c7573697a652c20343e005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243361646431376835666664656536393830656665666331450070616e69636b696e67006765745f756e636865636b65643c636f72653a3a666d743a3a72743a3a417267756d656e743e0064656275675f737472756374007b696d706c2332387d0065713c5b75385d2c205b75385d3e0044656275675475706c6500666d745f696e743c636f72653a3a666d743a3a6e756d3a3a55707065724865782c207536343e00636c616e67204c4c564d202872757374632076657273696f6e20312e37312e302d6e696768746c79202832663662633564323520323032332d30352d30392929006974657261746f72005f5a4e34636f726533737472313176616c69646174696f6e7331356e6578745f636f64655f706f696e74313768656364656330303032323838613566354500757466385f66697273745f627974650069735f636861725f626f756e64617279006d696e3c7573697a653e005f5a4e34636f72653373747235636f756e743330636f6e7461696e735f6e6f6e5f636f6e74696e756174696f6e5f627974653137686530636638653465356130663030393045005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137686134633765313364663063343439373145005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243361646431376833356564316564666234363437623138450077726974655f737472005f5a4e34636f726533666d74336e756d313247656e65726963526164697837666d745f696e743137686162643431393537653230363731373445006d617962655f756e696e697400696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e2c20636f72653a3a6f70733a3a72616e67653a3a52616e676546726f6d3c7573697a653e2c203132383e005f5a4e39395f244c5424636f72652e2e7374722e2e697465722e2e53706c6974496e636c7573697665244c54245024475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683536356238663563313134366339666645005f5a4e38315f244c5424636f72652e2e7374722e2e7061747465726e2e2e436861725365617263686572247532302461732475323024636f72652e2e7374722e2e7061747465726e2e2e53656172636865722447542431306e6578745f6d617463683137686231353436643361613035653433333145005f5a4e34636f72653463686172376d6574686f6473386c656e5f75746638313768343935363635353564666635366333654500656e636f64655f757466385f726177006172697468005f5a4e34345f244c54247538247532302461732475323024636f72652e2e6f70732e2e61726974682e2e52656d244754243372656d313768653539336133626230353330333763654500616c6c6f6300747261697473005f5a4e34636f726535736c6963653469746572313349746572244c54245424475424336e65773137683436326338393130346236666239373745005f5a4e34636f7265336e756d32335f244c5424696d706c24753230247573697a652447542431327772617070696e675f6d756c3137683933396664623563663661656266303945006e6577006d656d6368720077726170005f5a4e34636f726533666d74386275696c6465727331304465627567496e6e657235656e7472793137686361303935346134373764373230616545005f5a4e34636f726533666d74386275696c6465727331304465627567496e6e657235656e74727932385f24753762242475376224636c6f73757265247537642424753764243137686336663430636230393339663733626645005f5a4e34636f726533666d74336e756d313247656e65726963526164697837666d745f696e743137683330323730653937613764383866626145007061640070616e6963005f5a4e34636f726533666d74336e756d35335f244c5424696d706c2475323024636f72652e2e666d742e2e4c6f7765724865782475323024666f7224753230246936342447542433666d74313768663235653065383534373535336437314500696d7000616c7465726e617465006d6170005f5a4e3130325f244c5424636f72652e2e697465722e2e61646170746572732e2e6d61702e2e4d6170244c5424492443244624475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722447542434666f6c643137683439653563633739303661396231626645007772697465007b696d706c23377d006d696e5f62793c7573697a652c20666e28267573697a652c20267573697a6529202d3e20636f72653a3a636d703a3a4f72646572696e673e006765743c267374722c207573697a653e005f5a4e34636f726535736c69636535696e64657837345f244c5424696d706c2475323024636f72652e2e6f70732e2e696e6465782e2e496e646578244c542449244754242475323024666f72247532302424753562245424753564242447542435696e64657831376835623336343435386238326632343635450053706c6974496e7465726e616c006e6578743c636861723e0057726974650077726974655f636861723c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e007b696d706c2332367d005f5a4e34636f72653970616e69636b696e67313870616e69635f6e6f756e77696e645f666d743137683133386130386530383963323036303445005f5a4e34325f244c54242452462454247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d74313768633230363132656137383639386165344500666d74007b696d706c23307d004f7074696f6e007b696d706c23387d005f5a4e34636f726533707472376d75745f70747233315f244c5424696d706c2475323024244250246d757424753230245424475424336164643137686433383935323761353331303836366545006765745f756e636865636b65643c267374723e005f5a4e34636f726533666d7439466f726d6174746572313264656275675f73747275637431376838333134343030643138313466376534450070616e69635f737472005f5a4e34636f726533666d74386275696c64657273313564656275675f7475706c655f6e65773137683134383664383033383865636636373745005553495a455f4d41524b455200736c696365005f5a4e34636f7265336d656d377265706c6163653137683665313530623565366261663964346545007061645f696e74656772616c006765743c75383e005f5a4e34636f726535736c6963653469746572313349746572244c54245424475424336e65773137686231373834333338323430613463363745007b696d706c2331397d006e6578745f6d61746368005f5a4e34636f726536726573756c743139526573756c74244c542454244324452447542438616e645f7468656e3137686639613762303833656534636237383245005f5a4e37335f244c5424636f72652e2e666d742e2e6e756d2e2e5570706572486578247532302461732475323024636f72652e2e666d742e2e6e756d2e2e47656e657269635261646978244754243564696769743137683933663339316566393536306361643245005f5a4e34636f72653370747231303264726f705f696e5f706c616365244c542424524624636f72652e2e697465722e2e61646170746572732e2e636f706965642e2e436f70696564244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c542475382447542424475424244754243137683465633534623435323134663763393045005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683334323336653433336537396333623345006c74006368617273005f5a4e34636f72653373747232315f244c5424696d706c247532302473747224475424336765743137686361316261643162613538333362626645006765743c636f72653a3a6f70733a3a72616e67653a3a52616e6765546f3c7573697a653e3e00706f73745f696e635f73746172743c7573697a653e005f5a4e37355f244c54247573697a65247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c54242475356224542475356424244754242447542431336765745f756e636865636b65643137686630663432666234656339376261626145006164643c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e006d6574686f6473005f5a4e34636f726533666d74386275696c64657273313050616441646170746572347772617032385f24753762242475376224636c6f737572652475376424247537642431376862353032353031383864353564626337450063617061636974795f6f766572666c6f7700666d745f753634005f5a4e36385f244c5424636f72652e2e666d742e2e6275696c646572732e2e50616441646170746572247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f7374723137686539366438303337316562386433343445005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243361646431376836343831303738333031643161616237450049746572005f5a4e34636f72653373747232315f244c5424696d706c2475323024737472244754243563686172733137683635643537336338666664393434333645005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f723130616476616e63655f62793137683837343136383366376333383664636245006e6578745f636f64655f706f696e743c636f72653a3a736c6963653a3a697465723a3a497465723c75383e3e005f5a4e39335f244c5424636f72652e2e736c6963652e2e697465722e2e4368756e6b73244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137686264343939663734373230663065386245004f7264006164643c267374723e007b696d706c23367d00616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23357d3a3a656e7472793a3a7b636c6f737572655f656e7623307d3e004465627567536574005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f666d743137683565373464633863623261616161323645007b696d706c23327d005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542434697465723137686331616261316236653465646465623545005f5a4e34636f726533666d7439466f726d6174746572336e65773137686165623034366666366431666231663445005f5a4e34636f72653370747239636f6e73745f70747233335f244c5424696d706c247532302424425024636f6e7374247532302454244754243361646431376838353436653232346135313966363633450064656275675f7374727563745f6e657700746f5f7538005f5a4e34636f726533636d7035696d706c7336395f244c5424696d706c2475323024636f72652e2e636d702e2e5061727469616c4571244c54242452462442244754242475323024666f7224753230242452462441244754243265713137683436393566636435376362636161326145005f5a4e34636f726533666d743577726974653137683537653362636463656237646630393145006578706563745f6661696c6564006c656e5f6d69736d617463685f6661696c006f707300696e7472696e736963730073756d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e005f5a4e34636f7265336d656d377265706c61636531376838363534306363336630326138396663450069735f6e6f6e653c7573697a653e00697465723c5b7573697a653b20345d3e00696e746f5f697465723c5b7573697a653b20345d3e005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683366313636623661373436326234373945005f5a4e34636f726533666d7432727438417267756d656e7433666d74313768363232636537653835383430326338654500666d745f696e743c636f72653a3a666d743a3a6e756d3a3a4c6f7765724865782c207536343e00657175616c3c75382c2075383e005f5a4e34636f726535736c696365366d656d63687231326d656d6368725f6e616976653137686363623962373463393862393633336245006d656d6368725f6e6169766500616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23347d3a3a66696e6973683a3a7b636c6f737572655f656e7623307d3e005f5f616c6c6f635f6572726f725f68616e646c657200636f6e73745f707472005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f723373756d313768616537613566613764646461346162384500757466385f69735f636f6e745f62797465006e6578743c636f72653a3a666d743a3a72743a3a417267756d656e743e005f5a4e34636f726533666d74386275696c64657273313664656275675f7374727563745f6e65773137686135363836656238343531653037323245005f5a4e34636f72653970616e69636b696e67313370616e69635f646973706c6179313768663965353336303933393038663832624500656e64735f776974683c636861723e0065713c75382c2075383e007b696d706c23347d005f5a4e34636f726533737472313176616c69646174696f6e733137757466385f69735f636f6e745f6279746531376861396331376363326537313134623836450073706c69745f61745f756e636865636b65643c75383e0073706c69745f61743c75383e005f5a4e34636f72653373747235636f756e74313873756d5f62797465735f696e5f7573697a653137683733663965326535343130353136333245006e6578743c636f72653a3a666d743a3a72743a3a506c616365686f6c6465723e00417267756d656e74005f5a4e37355f244c54247573697a65247532302461732475323024636f72652e2e736c6963652e2e696e6465782e2e536c696365496e646578244c54242475356224542475356424244754242447542431336765745f756e636865636b6564313768656630633435353430343632353962624500636f6e7461696e735f7a65726f5f62797465005f5a4e37395f244c5424636f72652e2e726573756c742e2e526573756c74244c5424542443244524475424247532302461732475323024636f72652e2e6f70732e2e7472795f74726169742e2e54727924475424366272616e63683137683034646133323232663535363066313845005f5a4e34636f7265366f7074696f6e31336578706563745f6661696c65643137686332333330616533386638616564396545005f5a4e34636f726533707472376d75745f70747233315f244c5424696d706c2475323024244250246d7574247532302454244754243361646431376837336363316163653933303039363536450073756d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e2c207573697a653e005f5a4e35365f244c54247573697a65247532302461732475323024636f72652e2e697465722e2e7472616974732e2e616363756d2e2e53756d244754243373756d32385f24753762242475376224636c6f73757265247537642424753764243137683665653564323561643365666465373945007369676e5f61776172655f7a65726f5f70616400726561643c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e006e6578743c7573697a653e00756e777261705f6f723c267374723e005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243136616c69676e5f746f5f6f6666736574733137683265333033653231353164623038353745005f5a4e34636f726535736c69636532395f244c5424696d706c2475323024247535622454247535642424475424336765743137683037666466393631613031323632356145006e65773c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e007b696d706c2334347d0070616e69635f6e6f756e77696e645f666d740077726974655f7374723c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e577269746524475424313077726974655f636861723137683239666437616639333939643762333645005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243135636f70795f66726f6d5f736c69636531376c656e5f6d69736d617463685f6661696c3137686531663934356265353831313135613845006c6962726172792f616c6c6f632f7372632f6c69622e72732f402f616c6c6f632e643733613839653266303538366464312d6367752e30004974657261746f7200636f756e745f6368617273005f5a4e34636f72653469746572386164617074657273336d6170386d61705f666f6c6432385f24753762242475376224636c6f73757265247537642424753764243137686265643362346664336632356561633645005f5a4e34636f7265366f7074696f6e31354f7074696f6e244c542454244754243769735f6e6f6e653137683036303537623832613939663564313445005f5a4e34636f726535736c69636532395f244c5424696d706c247532302424753562245424753564242447542438616c69676e5f746f3137686361663565313535373365303734303345007b696d706c2331317d005f5a4e34636f726533636d70366d696e5f62793137683961363365346463336265666132393045005f5a4e34636f7265336d656d31326d617962655f756e696e697432304d61796265556e696e6974244c54245424475424357772697465313768643262633963366561386361383161624500656e636f64655f75746638005f5a4e34636f726533666d743557726974653977726974655f666d743137683364623431343565346436363932376245006669656c64007b696d706c2334307d005f5a4e36305f244c5424636f72652e2e63656c6c2e2e426f72726f774572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137686163386261333334363731373261333845005f5a4e34636f726533666d74336e756d35325f244c5424696d706c2475323024636f72652e2e666d742e2e4c6f7765724865782475323024666f72247532302469382447542433666d743137683039663834613031663936303437366145006e6578743c75383e00746f5f7573697a65006d656d005f5a4e34636f7265337074723577726974653137683934303032343231393363646338316545005f5a4e38395f244c5424636f72652e2e6f70732e2e72616e67652e2e52616e6765244c54245424475424247532302461732475323024636f72652e2e697465722e2e72616e67652e2e52616e67654974657261746f72496d706c2447542439737065635f6e65787431376834303038636235396134653064623339450061735f7573697a65006164643c636f72653a3a666d743a3a72743a3a417267756d656e743e00696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e005f5a4e34636f7265336e756d32335f244c5424696d706c24753230247573697a652447542431327772617070696e675f73756231376838643635306338643866353735643162450069735f70726574747900616461707465727300726561643c636861723e007b696d706c23337d00636861725f696e646963657300616c69676e5f746f3c75382c207573697a653e007772617070696e675f6d756c0077726974653c75383e005f5a4e35305f244c5424753634247532302461732475323024636f72652e2e666d742e2e6e756d2e2e446973706c6179496e742447542435746f5f75383137683636316463333963356464386666653545007061747465726e0069735f7375666669785f6f66005f5a4e34636f726535736c696365366d656d63687231346d656d6368725f616c69676e6564313768643864383232303663636532343531614500526573756c740050616441646170746572005f5a4e34636f726533666d7439466f726d6174746572337061643137683433336537613934646232626438653245005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f7374723137683865303931326361326264646233386345005f5a4e34636f726533666d7432727431325553495a455f4d41524b455232385f24753762242475376224636c6f7375726524753764242475376424313768643137376134333532613130653633314500466e4f6e6365006e756d005f5a4e38315f244c5424636f72652e2e7374722e2e697465722e2e4368617273247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f722447542435636f756e743137686638633866336432633063356164333545005f5a4e34636f726533666d7439466f726d617474657231397369676e5f61776172655f7a65726f5f7061643137683136323439616566366630343733333545006e65773c75383e007b696d706c23357d005f5a4e34636f726533636d70334f7264336d696e31376861623865636338303366663033636364450072756e005f5a4e34636f726533666d74386275696c64657273313044656275675475706c653969735f7072657474793137683131646663373739346165376162303045005f5a4e34636f726533666d7439466f726d617474657231327061645f696e74656772616c313277726974655f70726566697831376838346635386564303837613362643933450066756e6374696f6e00466f726d61747465720066696c746572006d61705f666f6c64005f5a4e38315f244c5424636f72652e2e7374722e2e697465722e2e4368617273247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683064323235303663643135633337363345007b696d706c2337307d005f5a4e39315f244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c54245424475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683634663237353939353136663335636545005f5a4e35355f244c542424524624737472247532302461732475323024636f72652e2e7374722e2e7061747465726e2e2e5061747465726e24475424313269735f7375666669785f6f663137686536396533336230613062663235373545007772617070696e675f7375620077726974655f666d743c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e005f5a4e35616c6c6f63377261775f766563313763617061636974795f6f766572666c6f7731376837363964333737343539393364316265450063616c6c5f6f6e63653c636f72653a3a666d743a3a72743a3a5553495a455f4d41524b45523a3a7b636c6f737572655f656e7623307d2c2028267573697a652c20266d757420636f72653a3a666d743a3a466f726d6174746572293e0062000000020000000000740000003400000063617061636974795f6f766572666c6f77002f0000007261775f76656300590000005f5f72646c5f6f6f6d004f000000616c6c6f6300540000005f5f616c6c6f635f6572726f725f68616e646c65720000000000f31b0000020074000000282600006a01000077726974653c636861723e00e22100006d617962655f756e696e697400bf2400006272616e63683c28292c20636f72653a3a666d743a3a4572726f723e00e90000006d75745f70747200c0220000696e736572743c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e00070400007b696d706c2334317d00ed1b0000636f70795f6e6f6e6f7665726c617070696e673c75383e005d060000466f726d617474657200ab2300007b696d706c2331377d00cc1f0000737065635f6e6578743c7573697a653e00701c0000706f73745f696e635f73746172743c7573697a653e00a71b0000617269746800d8180000446562756753657400091b00007b696d706c2332357d008d240000526573756c7400e72000006e6578745f636f64655f706f696e743c636f72653a3a736c6963653a3a697465723a3a497465723c75383e3e0034000000726561645f766f6c6174696c653c7573697a653e00151d0000697465723c5b7573697a653b20345d3e00d52100007265706c6163653c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e008d1f00007b636c6f7375726523307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e00e11c000073706c69745f61745f756e636865636b65643c75383e00c82100007265706c6163653c636861723e00a622000069735f6e6f6e653c7573697a653e002f1d00006765743c267374722c207573697a653e000d2500007b696d706c2332367d004321000069735f636861725f626f756e64617279006e240000726573756c7400581b000066756e6374696f6e00831f0000636f756e7400960600007061645f696e74656772616c00fb1c0000616c69676e5f746f5f6f6666736574733c75382c207573697a653e00751d00006c656e5f6d69736d617463685f6661696c00da0000006164643c75383e00581c00006e65773c75383e00fa030000646967697400211b0000666d743c28293e005523000070616e69636b696e6700b3220000756e777261705f6f723c267374723e0061200000636f6e7461696e735f6e6f6e5f636f6e74696e756174696f6e5f6279746500cd000000616c69676e5f6f66667365743c75383e00a71c00006e65773c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e000c2400007b696d706c2331397d00462300007772617070696e675f737562006f060000616c7465726e61746500322200006c74005a1f00006d61705f666f6c64006d20000073756d5f62797465735f696e5f7573697a6500ae010000417267756d656e7400e72100004d61796265556e696e6974009a050000666d7400b11b000072656d00ce2200006578706563745f6661696c656400f1020000666d745f696e743c636f72653a3a666d743a3a6e756d3a3a4c6f7765724865782c2075383e00bb1e0000636f6e7461696e735f7a65726f5f62797465004f13000072756e00c22000007b696d706c2334347d00882100007b696d706c2332387d003313000077726974655f707265666978005d1b0000466e4f6e636500da1d00006765743c267374723e005b000000636f6e73745f70747200b32100006e6578745f6d6174636800631d00006765743c75382c20636f72653a3a6f70733a3a72616e67653a3a52616e67653c7573697a653e3e00e5020000666d745f696e743c636f72653a3a666d743a3a6e756d3a3a55707065724865782c2075383e001322000077726974653c75383e00340100006164643c7573697a653e00471c00004974657200dd14000064656275675f7374727563745f6e6577001c1b00007b696d706c2335337d00b30000006164643c636f72653a3a666d743a3a72743a3a417267756d656e743e0009200000737472007323000070616e69635f646973706c61793c267374723e00ba1c0000697465723c75383e00701d0000636f70795f66726f6d5f736c69636500431f00006d617000832100007061747465726e00d9020000666d745f696e743c636f72653a3a666d743a3a6e756d3a3a4c6f7765724865782c207536343e005617000066696e69736800f50300007b696d706c2332397d00ac240000616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23347d3a3a66696e6973683a3a7b636c6f737572655f656e7623307d3e0073240000756e777261705f6661696c6564000a1c00006e6578743c75383e00af20000053706c6974496e7465726e616c003d200000646f5f636f756e745f6368617273003a1c00006e6578743c636f72653a3a666d743a3a72743a3a417267756d656e743e00fb1b0000736c696365006a17000044656275675475706c6500881f0000746f5f7573697a65004c1c0000706f73745f696e635f73746172743c75383e007a2000006974657200291f000073756d002d2200007b696d706c2335347d007d1c00007b696d706c2337307d00ce1d00006765745f756e636865636b65643c636f72653a3a666d743a3a72743a3a417267756d656e743e009f240000616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23357d3a3a656e7472793a3a7b636c6f737572655f656e7623307d3e00551a00007b696d706c23307d002b200000636861725f636f756e745f67656e6572616c5f6361736500a021000069735f7375666669785f6f66004d1f0000666f6c643c7573697a652c20636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c207573697a652c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e0025120000777261705f6275663c636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23317d3a3a777261703a3a7b636c6f737572655f656e7623307d3e00da1a000077726974655f666d743c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e00e3010000666d745f753634002a000000636f726500081d000061735f6368756e6b733c7573697a652c20343e000813000064656275675f7475706c655f6669656c64315f66696e697368009c0100005553495a455f4d41524b4552003e1f00006164617074657273002c2300007772617070696e675f6d756c002e1f00007b636c6f7375726523307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e004f2100006765743c636f72653a3a6f70733a3a72616e67653a3a52616e6765546f3c7573697a653e3e00a60000006164643c5b7573697a653b20345d3e00771f0000636f756e743c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e00951c0000696e746f5f697465723c5b7573697a653b20345d3e00dd1e0000666f6c643c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a6d61703a3a6d61705f666f6c643a3a7b636c6f737572655f656e7623307d3c2675382c207573697a652c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e3e00871800007b696d706c23317d008b23000070616e69635f6e6f756e77696e645f666d7400ed25000063686172006d1f000066696c746572009d1f0000656e756d657261746500971e00006d656d6368725f6e61697665008906000070616464696e67002e0300007b696d706c2336347d00181f00007b696d706c2334387d008c1800007772617000ca19000064656275675f7475706c655f6e657700e91400007b696d706c23327d00b301000061735f7573697a65001d1f000073756d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e0028220000696d706c7300ac1b00007b696d706c233232357d00131f0000616363756d00d81900005772697465005a23000070616e6963002e1c00006e6578743c636f72653a3a666d743a3a72743a3a506c616365686f6c6465723e0029210000636861727300531b00006f707300f22500006d6574686f647300781e000065713c75382c2075383e00c72000006e6578743c636861723e00950500007b696d706c2336357d005c210000656e64735f776974683c636861723e00c32100006d656d009b2100007b696d706c23337d007f23000070616e69635f737472007c1700006669656c64006e2200004f72640097010000727400de010000696d7000a71f00006e6578743c636f72653a3a736c6963653a3a697465723a3a497465723c636f72653a3a666d743a3a72743a3a506c616365686f6c6465723e3e00221c00006e6578743c7573697a653e00a21c0000497465724d75740069130000777269746500491d0000656e64735f776974683c75383e00b118000069735f70726574747900161c00006e6578743c5b7573697a653b20345d3e009f1800004465627567496e6e657200dd180000656e74727900f71e0000616476616e63655f62793c636f72653a3a7374723a3a697465723a3a43686172496e64696365733e00d402000047656e657269635261646978006a21000074726169747300fd020000666d745f696e743c636f72653a3a666d743a3a6e756d3a3a55707065724865782c207536343e005a1a000077726974655f7374723c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e00a22000006e65787400ea1e000073756d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e2c207573697a653e003e1700007b696d706c23347d00ee14000077726974655f73747200f72500006c656e5f75746638005222000065713c5b75385d2c205b75385d3e005d010000726561643c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e00ee1c000073706c69745f61743c75383e00b42000006e6578745f696e636c75736976653c636861723e001c0300007b696d706c2331317d0050010000726561643c636861723e007f090000706164005f1f00007b636c6f7375726523307d3c2675382c207573697a652c207573697a652c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e2c20636f72653a3a697465723a3a7472616974733a3a616363756d3a3a7b696d706c2334387d3a3a73756d3a3a7b636c6f737572655f656e7623307d3c636f72653a3a697465723a3a61646170746572733a3a6d61703a3a4d61703c636f72653a3a736c6963653a3a697465723a3a497465723c75383e2c20636f72653a3a697465723a3a61646170746572733a3a66696c7465723a3a7b696d706c23327d3a3a636f756e743a3a746f5f7573697a653a3a7b636c6f737572655f656e7623307d3c2675382c20636f72653a3a7374723a3a636f756e743a3a636861725f636f756e745f67656e6572616c5f636173653a3a7b636c6f737572655f656e7623307d3e3e3e3e00731a000077726974655f636861723c636f72653a3a666d743a3a6275696c646572733a3a506164416461707465723e00f3200000757466385f66697273745f6279746500bf1800007b696d706c23357d00b31f00006e6578743c636f72653a3a736c6963653a3a697465723a3a497465723c636f72653a3a666d743a3a72743a3a417267756d656e743e3e00612200006d696e5f62793c7573697a652c20666e28267573697a652c20267573697a6529202d3e20636f72653a3a636d703a3a4f72646572696e673e00ff1100006e657700152300006e756d007701000077726974653c636f72653a3a666d743a3a72743a3a416c69676e6d656e743e00b81d0000696e64657800942200004f7074696f6e009922000069735f736f6d653c7573697a653e00d81400006275696c646572730036210000636861725f696e646963657300a623000063656c6c00c00000006164643c267374723e00c71c00006765743c75382c207573697a653e00f31d00007b696d706c23367d00411e00006765743c75383e005b1700007b636c6f7375726523307d00db200000757466385f69735f636f6e745f6279746500d81e00004974657261746f7200621b000063616c6c5f6f6e63653c636f72653a3a666d743a3a72743a3a5553495a455f4d41524b45523a3a7b636c6f737572655f656e7623307d2c2028267573697a652c20266d757420636f72653a3a666d743a3a466f726d6174746572293e00a31e00006d656d6368725f616c69676e656400d41c0000616c69676e5f746f3c75382c207573697a653e00221d00006765745f756e636865636b65643c636f72653a3a666d743a3a72743a3a417267756d656e742c207573697a653e00410100006164643c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e00aa1d0000697465725f6d75743c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e008f2200006f7074696f6e0004260000656e636f64655f757466385f72617700d620000076616c69646174696f6e7300501e0000636d70007421000067657400e61d00006765745f756e636865636b65643c267374723e00291300007b696d706c23377d00051c00007b696d706c233138317d00d31e00006974657261746f72001812000064656275675f737472756374002f1e0000696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e2c20636f72653a3a6f70733a3a72616e67653a3a52616e676546726f6d3c7573697a653e3e00041f00006e74683c636f72653a3a7374723a3a697465723a3a43686172496e64696365733e0016260000656e636f64655f75746638007518000050616441646170746572008b1e00006d656d636872006f2100007b696d706c23387d00c11b0000696e7472696e7369637300ff240000696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e2c20636f72653a3a6f70733a3a72616e67653a3a52616e676546726f6d3c7573697a653e2c203132383e00c21f000072616e676500d32400007b696d706c2331357d007c0600007369676e5f61776172655f7a65726f5f70616400620600007369676e5f706c7573002f000000707472004100000064726f705f696e5f706c6163653c26636f72653a3a697465723a3a61646170746572733a3a636f706965643a3a436f706965643c636f72653a3a736c6963653a3a697465723a3a497465723c75383e3e3e001f200000636f756e745f636861727300641c00006e65773c5b7573697a653b20345d3e0016130000506f737450616464696e670017210000757466385f6163635f636f6e745f6279746500f81d0000696e6465783c636f72653a3a6d656d3a3a6d617962655f756e696e69743a3a4d61796265556e696e69743c75383e3e00402200007b696d706c23397d005c130000676574636f756e740092240000616e645f7468656e3c28292c20636f72653a3a666d743a3a4572726f722c2028292c20636f72653a3a666d743a3a6275696c646572733a3a7b696d706c23347d3a3a6669656c643a3a7b636c6f737572655f656e7623307d3e00812200006d696e3c7573697a653e0021030000746f5f753800ce0400007b696d706c2334307d005a1e0000657175616c3c75382c2075383e00ce240000617272617900000000000e00000002000000000074000000000000000e0000000200740000002826000000000000412a000000726973637600012000000004100572763634693270305f6d3270305f613270305f633270300084000000040040000000010101fb0e0d0001010101000000010000016c6962726172792f616c6c6f632f73726300007261775f7665632e727300010000616c6c6f632e72730001000000000902326e010000000000038a040105050a030109020001090c000001010402000902406e010000000000038d0301050d0a030b09020001090c00000101781e000004005e030000010101fb0e0d0001010101000000010000016c6962726172792f636f72652f7372632f6f7073006c6962726172792f636f72652f7372632f707472006c6962726172792f636f72652f7372632f666d74006c6962726172792f636f72652f737263006c6962726172792f636f72652f7372632f736c6963652f69746572006c6962726172792f636f72652f7372632f697465722f747261697473006c6962726172792f636f72652f7372632f737472006c6962726172792f636f72652f7372632f69746572006c6962726172792f636f72652f7372632f697465722f6164617074657273006c6962726172792f636f72652f7372632f6d656d006c6962726172792f636f72652f7372632f6d6163726f73006c6962726172792f636f72652f7372632f736c696365006c6962726172792f636f72652f7372632f6e756d006c6962726172792f636f72652f7372632f6172726179006c6962726172792f636f72652f7372632f63686172000066756e6374696f6e2e7273000100006d6f642e72730002000072742e7273000300006e756d2e727300030000636f6e73745f7074722e727300020000696e7472696e736963732e7273000400006d75745f7074722e7273000200006d6f642e7273000300006d6163726f732e7273000500006974657261746f722e72730006000076616c69646174696f6e732e727300070000616363756d2e727300060000636d702e72730004000072616e67652e7273000800006d61702e72730009000066696c7465722e727300090000636f756e742e727300070000697465722e7273000700006d6f642e7273000a00006f7074696f6e2e7273000400006d6f642e7273000b00006d6f642e727300070000696e6465782e7273000c00007472616974732e7273000700006d6f642e7273000c000075696e745f6d6163726f732e7273000d0000697465722e7273000c000070616e69636b696e672e727300040000656e756d65726174652e72730009000063656c6c2e7273000400006275696c646572732e727300030000726573756c742e7273000400006d617962655f756e696e69742e7273000a00006d6f642e7273000e0000636d702e7273000c00007061747465726e2e7273000700006d656d6368722e7273000c00006d6574686f64732e7273000f000061726974682e727300010000000009022ab301000000000003f90101040205090a03860a090000010403050503d3750902000109020000010104020009022eb301000000000003ea030105010a030009000001090200000101040400090230b301000000000003d2010105170a03130906000106039a7e0918000103e60109040001039a7e0924000105150603e80109020001051e0302090e00010405050d03b505091a00010406050903d20d090200010404051e03fa6c0904000104060509038613090400010405050d03ae72090800010406050903d20d090200010404051503fb6c09080001040605090385130902000106030009040001040405170603f56c0908000106039a7e0906000105140603f901090400010515030209040001051e037f091c000105150302090400010405050d03a305090200010406050903d20d090200010407050d039c73090c00010406050903e40c0902000106038f6b090a000104040514060381020902000105150301090400010407050d038b06090800010404051503f67909020001051e0302090a000105150301090200010405050d039905090400010406050903d20d090200010407050d039c73090c00010406050903e40c0902000106038f6b090800010407050d06038d08090400010404053e03827a09060001050d030209020001050a030109140001060b030009020001090400000101040800090272b401000000000003dd090105090a03e003091e0001051303a77c090c000106039b76090c000105090603f70d09040001051303ee7b0904000105190305090200010603967609020001050f0603fb0909020001050906030009020001038576090400010409051806038601090200010603fa7e09040001040a05150603b113090400010407050d03dc7409040001040b0505038c78090200010409051803ed0009080001040c051c03af7f090200010409051803d100090200010408050d03e50809020001050f031009020001050906030009020001052306030909020001051a06030009040001050906038d0409040001051a03f97b09020001051b03e90009020001053103a47f09060001051503dc000904000106038d7509060001050606039d0a09200001060b0300091c0001050003e3750904000104020509060394090926000106030009060001040805110603f900090400010402050903cd00090a000106030009040001040805110603b37f090400010603f3750914000105090603800b09020001040d05340353090600010408050d032e090400010603ff740910000105150603f30a090200010530030a0904000105230603000904000105300300090200010383750906000105090603800b090c0001040d0534035309040001040e050c039a7a090200010408050d039406090200010603ff74090c000105240603970a090a00010511030109040001030109140001050903fb7e090e0001040d053403bf01090800010408050d03c27e09080001051103fa00091000010603f175091000010603910a090200010301090400010603ee7509080001040d05340603d30a09020001090600000101040800090256b601000000000003f2090105140a0301091c0001051103010904000105140302090e0001052c060300090200010b03000912000103897609040001050a0603f80909020001060b0300090a00010904000001010408000902acb601000000000003bb0a01041405120a039b7a090200010408050c03e7050916000104150509039a78090200010408050c03e607090800010518030509040001051d060300090400010405050d0603dc7c09040001040a050903b87b09040001040b05000603a97d09120001041205260603910109040001051106030009020001040a05100603c70109040001040d053403fb0709040001040e050c039a7a090200010409051803997c09020001040b050d03a07f0904000105080301090800010516030a090400010505035b0904000105110306090400010508032109040001051a0305090400010505035a090400010511060300090200010505030009040001050c06032909040001051e030509040001051203010904000105050351090400010511060300090200010505030009040001050d06032f090400010412050903cb00090200010603f47e090400010409051806038601091e0001040b050d03a07f090400010508030109040001060359090400010603330908000106034d09040001050c06033b09040001050006034509040001051a060338090400010511035a0904000106030009040001051e06032e09040001051203010904000105050351090400010511060300090600010505030009040001050d06032f090200010412050903cb00090600010416050c03cc000904000105090304090200010417050c037d0904000104160513030f0904000104180509032c090800010603ec7d0904000104140603bc0709020001041803d87a090400010603ec7d0904000104140603bc07090200010603c4780902000104080603d40a0904000105120304090400010411050803c37509080001060365090400010409051806038601090200010603fa7e09040001040a05150603b113090400010407050d03dc7409040001040b0505038c78090200010409051803ed0009080001040c051c03af7f090200010409051803d100090200010402051f03bb0c0904000104190545036509060001051603800e090800010409051803e065090600010603fa7e09040001040a05150603b113090200010407050d03dc7409040001040b0505038c78090200010409051803ed0009080001040c051c03af7f090200010409051803d100090200010603fa7e090200010386010902000103fa7e09020001040a05150603b113090600010407050d03dc7409040001040b0505038c78090200010409051803ed0009080001040c051c03af7f090200010409051803d100090200010603fa7e09020001041105150603c7000922000105000603b97f09060001051b0603fe00090e00010534060300090400010533030009020001051b030009040001041a050d0603e7080902000104110505039a77090400010509035b09020001050c030609020001041b03e80a090200010603b874090200010419053806039908091200010405050d03867f090400010409051803e779090600010603fa7e09020001041105190603d0000904000105120301090200010507032309020001050606030009040001051203000902000106035d09020001050503230902000105110360090400010507032009020001050606030009040001051206035d090200010323090200010505060300090200010507030009040001050603000904000105120300090200010505030009020001051206035d0902000105050323090200010511036009020001050703200904000105060603000904000105120300090200010505030009020001040905180603120904000104110511034e09040001040905180332090200010603000906000103fa7e090400010386010904000103fa7e09040001038601090600010411051206035d090600010407050d03aa07090200010411050703e7780902000105060603000904000105120300090200010505030009020001040905180603120904000104110511035e09020001040905180322090200010603fa7e090400010411051b0603fe00090200010534060300090400010533030009020001051b030009040001041a050d0603e7080902000104110505039a7709040001050d0367090200010408051403f60909020001051b0317090400010535037009060001051503100904000106038d750906000103f30a09260001053006030a0904000105230603000904000105300300090200010383750906000105090603800b090e0001040d0534035309040001040e050c039a7a090200010408050d039406090200010603ff74090c000105280603e30a090a00010515030109040001050903b07e090e0001040d053403bf0109080001040e050c039a7a090400010408050d03a804090400010603eb7609100001040d05340603d30a0902000104080506031609040001060b030009140001090400000101041c00090224ba01000000000003ed000105050a030709020001090c00000101040800090232ba01000000000003b7080105090a03bb7909180001050b03c90609080001050903b77909040001050503c90609080001050e030e090200010409051803bc78090400010603fa7e0904000103860109040001040805150603cb0709220001051406030009020001051506030109020001052d0603000904000105150300090400010510060313090600010505060300090200010511060301090200010505060300090400010511060301090400010533036f09020001050503110904000105150304090200010505030f090600010403050c039978090600010603ed7e090a0001051d0603960109040001051b0603000902000103ea7e09020001040805090603eb080902000105190301090400010505030e090800010403050c039978090600010603ed7e090a0001051d0603960109040001051b0603000902000103ea7e09020001040805090603ec0809020001052d0307090400010405050d03ac7e090200010403050903eb7909040001051a060300090200010509030009020001040805110603cc07090400010409051803b078090200010408051d03b907091000010409051803c778090400010603fa7e0904000103860109080001040805150603bd0709120001051406030009020001051506030109020001052d060300090400010515030009040001040305090603c67809060001051a060300090200010509030009040001040805110603bc07090400010409051803c078090200010408051a03d707090a00010417050c03fc78090400010603a77e090600010408051a0603dd08090200010417050c03fc78090400010408051a038407090400010405050d03c27e090400010408050903bf0109040001052106030009040001050903000908000103a2770906000105020603e20809060001060b030009100001090400000101041e000902b0bb01000000000003ba0501040805090a03ba0609000001091200000101041e000902c2bb01000000000003d50501040805090a039f06090000010912000001010420000902d4bb01000000000003f10c0105050a030109020001090c000001010414000902e2bb010000000000038a0f01041c05050a038b7209020001090c00000101041c000902f0bb01000000000003cf0001050e0a031009020001090c000001010404000902febb010000000000039901010407050d0a03f30609060001040405000603f3770908000106039301090800010421050903d602090200010404051403ea7c090400010603ad7f09080001052306032a0902000103e900090800010603ed7e090400010417050c0603ed03090a00010404050903817d090a0001050e032e09160001060b0300090200010417050d0603d20209040001090e00000101041f0009026ebc010000000000031e010412050c0a03ce040946000104190523039c0d091800010423050d03d26e09040001041f034a090a00010301090400010412050c03c704090e00010424051903b17e090800010417050c0342090a00010425050803cb7d09080001050b030d0906000106034809040001050c0603390902000105090304090c0001050b037b090200010402051f03890d09060001051b03010908000104250508039273090400010603ac7f090e000105100603eb00090600010405050d03b406090400010425051503c679090400010529030409060001041a050d03e508090200010425050503c67609020001051503d2000908000105290304090a0001041a050d03e408090200010425050503c67609020001050903db0009080001050b037209020001050c03580906000105090304090c0001050b037b09020001060348090400010603e1000904000106039f7f09040001050c06033909060001050b037f090c000106034809080001042405200603b403090200010511060300090200010417050c0603ac7f090800010423050d03fb7d090200010424051c03dd02090400010603c87c09040001041f051006032109140001051103010906000106035e090e00010419050906038912090800010603f76d09040001041f050606032a09100001060b0300091a000109040000010104080009022abe01000000000003a20101052b0a0301090c00010426050803f60b09020001050d031f09040001050f0363090800010513032009060001050d06030009040001051206030109080001050d06030009040001050f060361090c00010513032209060001050d06030009040001051206030109080001050d06030009060001051206030109080001050d060300090400010512060303090c0001050d06030009060001051206030109080001050d06030009060001051206030109080001050d06030009060001051206030109080001050d06030009040001040805090603dc73090a000105060301090a0001060b0300090200010904000001010408000902debe01000000000003be010105090a0301090200010506030109300001060b030009020001090400000101040800090216bf01000000000003c5010105090a030109000001090a00000101040800090220bf01000000000003c9010105090a030109020001052b0359090c00010426050803f60b09020001050d031f09040001050f0363090800010513032009060001050d06030009040001051206030109080001050d06030009040001050f060361090c00010513032209060001050d06030009040001051206030109080001050d06030009060001051206030109080001050d060300090400010512060303090c0001050d06030009060001051206030109080001050d06030009060001051206030109080001050d06030009060001051206030109080001050d06030009040001040805090603dc73090a000105060328090a0001060b0300090200010904000001010408000902d6bf01000000000003cd010105090a0301090200010371091e00010506031009140001060b030009020001090400000101041f00090210c001000000000003b3020105170a0301091200010420050903f10709040001041f03a078090200010603ba7d0908000105100603b602090400010408050903c10b09040001041f050006038972090400010408050903f70d09040001041f05100603bf740904000105000603ca7d09020001051e0603c002090400010603c07d0904000105140603b702090a00010408050903be0909040001041f051503c376091600010603c87d09020001040805090603f50b090e0001041f051e03cb76090a00010408050903b50909020001042003a70309040001041f051103a673090200010408051403e406090c00010603da7609040001041f05210603bb02090200010408051703e806090400010414050903f002090800010408051303947d090a0001051403010904000103010904000105180301090800010509037709080001041f0511039c79091400010408050903e40609040001041f0511039c79090a00010408050903b80909080001041f050006038b740912000105090603b502090200010311090400010506030209060001060b030009100001090400000101041f00090230c101000000000003d3030105170a03a87f091200010420050903aa0709080001041f03d67809020001031209040001050603c90009040001060b03000910000103a97c0904000105100603fd02090400010408050903fa0a09040001041f050006038972090400010408050903f70d09040001041f051006038675090400010514030a090200010408050903ee0809020001041f051503937709180001051103020902000105140374090a00010408050903f70809020001041f0515038a77091800010408051403a706090200010603da7609040001041f052106038203090200010408051703a106090400010414050903f002090800010408051303947d090a0001051403010904000103010904000105180301090800010509037709080001041f051103e379091e00010408050903f10809080001091600000101040800090230c201000000000003e40f0105090a03907c090c0001041f050503a376090c00010408050903cf0d090c0001041f050c03fd72090e0001050006039c7d09020001050c03e40209040001039c7d09020001042005090603a60a09020001041f051403c07809020001050006039a7d090a0001051403e60209020001040805090603910b09080001041f051403ef740906000104080509038f0909020001041f051503f2760914000104080509038e0909020001041f03f776091600010408050603fd0c09040001060b0300090a00010904000001010419000902c8c2010000000000038a1a01050d0a030109020001090c000001010404000902d6c2010000000000039901010407050d0a03f30609060001040405000603f3770908000106039401090c00010421050903d502090200010404051403ea7c090400010427052d03ef03090800010404052303d27c090800010603ec7e090400010417050c0603ed03090a00010404050903817d090a0001050e032e09160001060b0300090200010417050d0603d20209040001090e00000101040400090248c3010000000000039901010407050d0a03f30609060001040405000603f3770908000106039301090c00010421050903d602090200010404051403ea7c090400010427052d03ef03090800010404052303d17c090800010603ed7e090400010417050c0603ed03090a00010404050903817d090a0001050e032e09160001060b0300090200010417050d0603d20209040001090e000001010408000902bac301000000000003cf110105090a03ec01090000010916000001010422000902d0c301000000000003820101040805090a03f20a090a00010422051e038f75090200010408050903f10a09020001041f050503a376091000010408050903cf0d090c0001041f050c03fd7209140001050006039c7d09020001050c03e40209040001039c7d09020001042005090603a60a09020001041f051403c07809020001050006039a7d090a0001051403e60209020001040805090603910b09080001041f051403ef740906000104080509038f0909020001041f051503f2760914000104080509038e0909020001041f03f776091600010422050f03977e09040001060b030009080001090400000101040400090272c4010000000000039901010407050d0a03f30609060001040405000603f3770908000106039401090800010421050903d502090200010404051403ea7c090400010603ad7f09080001052306032a0902000103ea00090800010603ec7e090400010417050c0603ed03090a00010404050903817d090a0001050e032e09160001060b0300090200010417050d0603d20209040001090e00000101004743433a2028292031322e322e30004c696e6b65723a204c4c442031362e302e320000000000000000000000000000000000000000000000000000000000000000010000000400f1ff00000000000000000000000000000000220000000000050038c902000000000000000000000000002b000000020004008a36010000000000640000000000000000000000000004008a36010000000000000000000000000000000000000004008c360100000000000000000000000000000000000000040094360100000000000000000000000000fc00000000000400a0360100000000000000000000000000080100000200040086c801000000000056000000000000006701000002000400106e01000000000008000000000000000000000000000400ee3601000000000000000000000000007601000002000400ee3601000000000010000000000000000000000000000400ee3601000000000000000000000000000000000000000400fe360100000000000000000000000000c701000002000400fe36010000000000ee000000000000000000000000000400fe36010000000000000000000000000000000000000004000037010000000000000000000000000000000000000004000a3701000000000000000000000000004202000000000400d63701000000000000000000000000004e02000001000100e2090100000000002b00000000000000780200000200040024ba0100000000000e000000000000000000000000000400ec370100000000000000000000000000a502000002000400ec37010000000000d4040000000000000000000000000400ec3701000000000000000000000000000000000000000400ee370100000000000000000000000000000000000000040008380100000000000000000000000000f8020000020004001a47010000000000c600000000000000ce03000002000400043e01000000000030000000000000001f04000002000400343e01000000000030000000000000007404000002000400283d010000000000dc000000000000008f05000000000400563c01000000000000000000000000009b05000001000100690b0100000000003500000000000000c605000000000400643c0100000000000000000000000000d205000001000100410b0100000000002800000000000000fd05000002000400c8c20100000000000e0000000000000063060000000004007a3c01000000000000000000000000006f06000000000400903c01000000000000000000000000007b060000000004009e3c01000000000000000000000000008706000000000400a83c01000000000000000000000000009306000001000100f00a0100000000003000000000000000be06000000000400b63c01000000000000000000000000000000000000000400c03c0100000000000000000000000000ca06000002000400c03c01000000000068000000000000000000000000000400c03c01000000000000000000000000009207000002000400f0bb0100000000000e000000000000000000000000000400283d01000000000000000000000000000000000000000400283d010000000000000000000000000000000000000004002a3d01000000000000000000000000000000000000000400403d01000000000000000000000000000000000000000400043e01000000000000000000000000000000000000000400043e01000000000000000000000000000000000000000400063e01000000000000000000000000000000000000000400083e0100000000000000000000000000cd07000002000400086e0100000000000800000000000000da07000002000400286e0100000000000a000000000000000000000000000400343e01000000000000000000000000000000000000000400343e01000000000000000000000000000000000000000400363e01000000000000000000000000000000000000000400383e01000000000000000000000000000000000000000400643e0100000000000000000000000000f507000002000400643e0100000000007a010000000000000000000000000400643e01000000000000000000000000000000000000000400663e010000000000000000000000000000000000000004007e3e01000000000000000000000000005b08000000000400a23f01000000000000000000000000006708000001000100b90b01000000000033000000000000009208000000000400b03f01000000000000000000000000009f08000001000100ec0b0100000000002700000000000000ca08000000000400be3f0100000000000000000000000000d708000000000400c83f0100000000000000000000000000e408000001000100130c01000000000028000000000000000000000000000400de3f01000000000000000000000000000f09000002000400de3f010000000000aa010000000000000000000000000400de3f01000000000000000000000000000000000000000400e03f01000000000000000000000000000000000000000400fa3f010000000000000000000000000076090000000004005041010000000000000000000000000083090000010001003b0c0100000000003200000000000000ae090000000004005e410100000000000000000000000000bb090000010001006d0c0100000000002800000000000000e60900000000040068410100000000000000000000000000f30900000000040072410100000000000000000000000000000000000000040088410100000000000000000000000000000a0000020004008841010000000000c00100000000000000000000000004008841010000000000000000000000000000000000000004008a4101000000000000000000000000000000000000000400a4410100000000000000000000000000700a000000000400244301000000000000000000000000007d0a000001000100950c0100000000009100000000000000a80a00000000040032430100000000000000000000000000b50a000001000100260d0100000000002a00000000000000000000000000040048430100000000000000000000000000e00a0000020004004843010000000000820100000000000000000000000004004843010000000000000000000000000000000000000004004a4301000000000000000000000000000000000000000400644301000000000000000000000000003e0b000000000400b44401000000000000000000000000000000000000000400ca4401000000000000000000000000004b0b000002000400ca4401000000000050020000000000000000000000000400ca4401000000000000000000000000000000000000000400cc4401000000000000000000000000000000000000000400e644010000000000000000000000000000000000000004001a47010000000000000000000000000000000000000004001a47010000000000000000000000000000000000000004001c4701000000000000000000000000000000000000000400344701000000000000000000000000000000000000000400e04701000000000000000000000000000000000000000400e04701000000000000000000000000000000000000000400e447010000000000000000000000000000000000000004001848010000000000000000000000000000000000000004001848010000000000000000000000000000000000000004001a480100000000000000000000000000990c0000000004001a480100000000000000000000000000a60c00000100060088ca0200000000001000000000000000cf0c0000020004002cae010000000000c204000000000000080d00000200040006b301000000000024000000000000003f0d0000020004004c380200000000001c00000000000000b20d0000020004006838020000000000da00000000000000e80d0000020004007ac60100000000004e00000000000000300e000002000400204a0200000000008601000000000000710e0000020004004aac0100000000008200000000000000b20e000002000400243802000000000028000000000000002b0f000000000400824f0100000000000000000000000000380f0000010001000c050100000000001100000000000000640f000000000400c84f0100000000000000000000000000710f00000200040010aa010000000000c001000000000000a90f00000000040022500100000000000000000000000000b60f00000200040060930100000000007c00000000000000f80f000000000400ee5001000000000000000000000000000510000002000400daa901000000000036000000000000005f100000000004009a5101000000000000000000000000006c10000000000400d851010000000000000000000000000079100000000004000452010000000000000000000000000086100000000004001e5201000000000000000000000000009310000001000100d00401000000000021000000000000009c10000002000400faa30100000000002200000000000000171100000200040088a1010000000000d600000000000000ab110000020004001ca40100000000003a00000000000000e41100000200040052a501000000000042000000000000002312000000000400b25201000000000000000000000000003012000000000400ca5201000000000000000000000000003d12000001000100b0050100000000001c000000000000004712000000000400f0520100000000000000000000000000541200000200040056a4010000000000fc00000000000000dc120000020004008ea30100000000006c000000000000000f1300000200040058a6010000000000640000000000000062130000020004000e5002000000000054020000000000009a1300000200040058720100000000005800000000000000fa13000002000400fc4d0200000000009a000000000000002c140000020004005e7001000000000058000000000000008314000002000400ae6f0100000000005800000000000000df1400000200040006700100000000005800000000000000391500000200040042390200000000002a020000000000006e15000002000400fe6e0100000000005800000000000000cb15000002000400566f01000000000058000000000000002616000002000400b670010000000000580000000000000081160000020004004e6e0100000000005800000000000000dc16000002000400a66e01000000000058000000000000003517000002000400d4a801000000000072000000000000008b170000020004005ccf010000000000ba000000000000000c180000020004000e71010000000000520000000000000065180000020004009e3b02000000000018030000000000009c18000002000400da730100000000004e00000000000000fd180000020004000873010000000000860000000000000049190000020004008e730100000000004c000000000000009519000002000400b0720100000000005800000000000000e01900000200040060710100000000005800000000000000331a00000200040028740100000000009400000000000000941a000002000400d4590200000000007400000000000000c21a000002000400485a0200000000004a3a000000000000f61a000002000400d2450200000000004e04000000000000321b000002000400b8710100000000005200000000000000921b000002000400b63e0200000000008c03000000000000d61b0000020004000a720100000000004e00000000000000291c0000020004006ed1010000000000c000000000000000b51c00000200040062520200000000007207000000000000f41c000002000400424202000000000090030000000000003b1d000002000400964e0200000000007801000000000000701d000002000400bc740100000000009400000000000000d11d000000000400ba6c0100000000000000000000000000de1d000000000400ca6c0100000000000000000000000000eb1d00000100010000020100000000001c00000000000000f11d000000000400d66c0100000000000000000000000000fe1d0000010001005e0a0100000000002b00000000000000291e000000000400de6c0100000000000000000000000000361e00000100010040020100000000002000000000000000601e000002000400d4bb0100000000000e00000000000000931e000000000400f66c0100000000000000000000000000a01e000000000400026d0100000000000000000000000000ad1e000000000400146d0100000000000000000000000000ba1e0000000004001c6d0100000000000000000000000000c71e00000100010020020100000000002000000000000000f11e0000000004002e6d0100000000000000000000000000fe1e000000000400366d01000000000000000000000000000b1f000000000400406d0100000000000000000000000000181f000000000400486d0100000000000000000000000000251f000000000400526d0100000000000000000000000000321f0000000004005a6d01000000000000000000000000003f1f000000000400646d01000000000000000000000000004c1f000001000100200b01000000000021000000000000000000000000000400706d0100000000000000000000000000771f000002000400706d0100000000000a000000000000000000000000000400706d0100000000000000000000000000891f000002000400eeb2010000000000180000000000000000000000000004007a6d0100000000000000000000000000be1f0000020004007a6d010000000000080000000000000000000000000004007a6d0100000000000000000000000000c91f000002000400c299010000000000d4030000000000000000000000000400826d01000000000000000000000000005420000002000400826d01000000000008000000000000000000000000000400826d01000000000000000000000000006120000002000400969d010000000000f20300000000000000000000000004008a6d0100000000000000000000000000ee200000020004008a6d0100000000004e0000000000000000000000000004008a6d010000000000000000000000000000000000000004008c6d01000000000000000000000000000000000000000400966d01000000000000000000000000000000000000000400d86d0100000000000000000000000000fb20000002000400d86d01000000000030000000000000000000000000000400d86d01000000000000000000000000000000000000000400da6d01000000000000000000000000000000000000000400e06d01000000000000000000000000000000000000000400086e01000000000000000000000000000000000000000400086e01000000000000000000000000000000000000000400106e01000000000000000000000000000000000000000400106e01000000000000000000000000000000000000000400186e01000000000000000000000000000d21000002000400186e01000000000008000000000000000000000000000400186e01000000000000000000000000000000000000000400206e01000000000000000000000000001c21000002000400206e01000000000008000000000000000000000000000400206e01000000000000000000000000000000000000000400286e01000000000000000000000000000000000000000400286e01000000000000000000000000003021000002000400406e0100000000000e000000000000000000000000000400326e01000000000000000000000000003a21000002000400326e0100000000000e000000000000000000000000000400326e01000000000000000000000000000000000000000400326e01000000000000000000000000000000000000000400326e01000000000000000000000000000000000000000400346e01000000000000000000000000000000000000000400346e01000000000000000000000000000000000000000400366e01000000000000000000000000000000000000000400406e01000000000000000000000000000000000000000400406e01000000000000000000000000000000000000000400406e01000000000000000000000000000000000000000400406e01000000000000000000000000000000000000000400406e01000000000000000000000000000000000000000400426e01000000000000000000000000000000000000000400426e01000000000000000000000000000000000000000400446e010000000000000000000000000000000000000004004e6e010000000000000000000000000000000000000004004e6e010000000000000000000000000000000000000004004e6e01000000000000000000000000000000000000000400506e01000000000000000000000000000000000000000400546e0100000000000000000000000000732100000200040080cb0100000000006601000000000000ba2100000200040040ce010000000000a2000000000000005722000000000400866e010000000000000000000000000064220000000004008e6e01000000000000000000000000007122000001000100600201000000000020000000000000000000000000000400a66e01000000000000000000000000000000000000000400a66e01000000000000000000000000000000000000000400a86e01000000000000000000000000000000000000000400ac6e01000000000000000000000000009c22000000000400de6e0100000000000000000000000000a922000000000400e66e01000000000000000000000000000000000000000400fe6e01000000000000000000000000000000000000000400fe6e01000000000000000000000000000000000000000400006f01000000000000000000000000000000000000000400046f0100000000000000000000000000b622000000000400366f0100000000000000000000000000c3220000000004003e6f01000000000000000000000000000000000000000400566f01000000000000000000000000000000000000000400566f01000000000000000000000000000000000000000400586f010000000000000000000000000000000000000004005c6f0100000000000000000000000000d0220000000004008e6f0100000000000000000000000000dd22000000000400966f01000000000000000000000000000000000000000400ae6f01000000000000000000000000000000000000000400ae6f01000000000000000000000000000000000000000400b06f01000000000000000000000000000000000000000400b46f0100000000000000000000000000ea22000000000400e66f0100000000000000000000000000f722000000000400ee6f010000000000000000000000000000000000000004000670010000000000000000000000000000000000000004000670010000000000000000000000000000000000000004000870010000000000000000000000000000000000000004000c70010000000000000000000000000004230000000004003e70010000000000000000000000000011230000000004004670010000000000000000000000000000000000000004005e70010000000000000000000000000000000000000004005e7001000000000000000000000000000000000000000400607001000000000000000000000000000000000000000400647001000000000000000000000000001e23000000000400967001000000000000000000000000002b230000000004009e7001000000000000000000000000000000000000000400b67001000000000000000000000000000000000000000400b67001000000000000000000000000000000000000000400b87001000000000000000000000000000000000000000400bc7001000000000000000000000000003823000000000400ee7001000000000000000000000000004523000000000400f670010000000000000000000000000000000000000004000e71010000000000000000000000000000000000000004000e7101000000000000000000000000000000000000000400107101000000000000000000000000000000000000000400127101000000000000000000000000005223000002000400c2cd0100000000007e00000000000000d72300000000040040710100000000000000000000000000e42300000000040048710100000000000000000000000000000000000000040060710100000000000000000000000000000000000000040060710100000000000000000000000000000000000000040062710100000000000000000000000000000000000000040066710100000000000000000000000000f12300000000040098710100000000000000000000000000fe23000000000400a07101000000000000000000000000000000000000000400b87101000000000000000000000000000000000000000400b87101000000000000000000000000000000000000000400ba7101000000000000000000000000000000000000000400bc7101000000000000000000000000000b240000020004004acd01000000000078000000000000009124000000000400ea7101000000000000000000000000009e24000000000400f271010000000000000000000000000000000000000004000a72010000000000000000000000000000000000000004000a72010000000000000000000000000000000000000004000c720100000000000000000000000000000000000000040010720100000000000000000000000000ab2400000000040036720100000000000000000000000000b8240000000004003e72010000000000000000000000000000000000000004005872010000000000000000000000000000000000000004005872010000000000000000000000000000000000000004005a72010000000000000000000000000000000000000004005e720100000000000000000000000000c52400000000040090720100000000000000000000000000d224000000000400987201000000000000000000000000000000000000000400b07201000000000000000000000000000000000000000400b07201000000000000000000000000000000000000000400b27201000000000000000000000000000000000000000400b6720100000000000000000000000000df24000000000400e8720100000000000000000000000000ec24000000000400f072010000000000000000000000000000000000000004000873010000000000000000000000000000000000000004000873010000000000000000000000000000000000000004000a730100000000000000000000000000000000000000040010730100000000000000000000000000f92400000200040086ca0100000000006200000000000000322500000200040050cb010000000000300000000000000072250000000004006e7301000000000000000000000000007f250000000004007873010000000000000000000000000000000000000004008e73010000000000000000000000000000000000000004008e7301000000000000000000000000000000000000000400907301000000000000000000000000000000000000000400947301000000000000000000000000008c25000000000400b87301000000000000000000000000009925000000000400c07301000000000000000000000000000000000000000400da7301000000000000000000000000000000000000000400da7301000000000000000000000000000000000000000400dc7301000000000000000000000000000000000000000400e0730100000000000000000000000000a62500000000040006740100000000000000000000000000b3250000000004000e74010000000000000000000000000000000000000004002874010000000000000000000000000000000000000004002874010000000000000000000000000000000000000004002a74010000000000000000000000000000000000000004002e740100000000000000000000000000c025000002000400e6cc010000000000640000000000000005260000000004008474010000000000000000000000000012260000000004008c7401000000000000000000000000001f260000000004009c7401000000000000000000000000002c26000000000400a47401000000000000000000000000000000000000000400bc7401000000000000000000000000000000000000000400bc7401000000000000000000000000000000000000000400be7401000000000000000000000000000000000000000400c27401000000000000000000000000003926000000000400187501000000000000000000000000004626000000000400207501000000000000000000000000005326000000000400307501000000000000000000000000006026000000000400387501000000000000000000000000000000000000000400507501000000000000000000000000006d260000020004005075010000000000bc0000000000000000000000000004005075010000000000000000000000000000000000000004005275010000000000000000000000000000000000000004005a750100000000000000000000000000b0260000020004000c760100000000009a00000000000000f626000002000400a676010000000000dc0000000000000000000000000004000c76010000000000000000000000000000000000000004000c76010000000000000000000000000000000000000004000e76010000000000000000000000000000000000000004001676010000000000000000000000000038270000000004002c7601000000000000000000000000004527000001000100a00201000000000040000000000000000000000000000400a67601000000000000000000000000000000000000000400a67601000000000000000000000000000000000000000400aa7601000000000000000000000000000000000000000400b676010000000000000000000000000083270000020004008277010000000000ee1a000000000000000000000000040082770100000000000000000000000000c72700000000050040c90200000000000000000000000000d12700000000050048c90200000000000000000000000000db2700000000050050c90200000000000000000000000000e52700000000050058c90200000000000000000000000000ef2700000000050060c90200000000000000000000000000f92700000000050068c90200000000000000000000000000032800000000050070c902000000000000000000000000000d2800000000050078c9020000000000000000000000000000000000000004008277010000000000000000000000000000000000000004008477010000000000000000000000000000000000000004009e77010000000000000000000000000017280000000004001e78010000000000000000000000000024280000000004003278010000000000000000000000000031280000000004007e7801000000000000000000000000003e28000000000400927801000000000000000000000000004b28000000000400dc7801000000000000000000000000005828000000000400f678010000000000000000000000000065280000000004003c7901000000000000000000000000007228000000000400527901000000000000000000000000000000000000000400709201000000000000000000000000007f280000020004007092010000000000f00000000000000000000000000004007092010000000000000000000000000000000000000004007292010000000000000000000000000000000000000004007a9201000000000000000000000000000000000000000400609301000000000000000000000000000000000000000400609301000000000000000000000000000000000000000400629301000000000000000000000000000000000000000400689301000000000000000000000000000000000000000400dc930100000000000000000000000000bd28000002000400dc9301000000000014040000000000000000000000000400dc9301000000000000000000000000000000000000000400de9301000000000000000000000000000000000000000400f8930100000000000000000000000000ff28000002000400f0970100000000003c000000000000003929000000000400be9401000000000000000000000000004729000001000100c0030100000000001c00000000000000502900000200040036980100000000004c00000000000000892900000200040082980100000000004c00000000000000d429000002000400e2bb0100000000000e00000000000000072a00000000040036970100000000000000000000000000152a0000000004004a970100000000000000000000000000232a00000000040054970100000000000000000000000000312a0000000004005e9701000000000000000000000000003e2a000000000400689701000000000000000000000000004c2a00000100010060030100000000002100000000000000552a00000000040072970100000000000000000000000000632a000001000100900301000000000024000000000000006c2a000000000400809701000000000000000000000000007a2a0000000004008a970100000000000000000000000000882a00000100010030030100000000002100000000000000912a000000000400949701000000000000000000000000009f2a0000000004009e970100000000000000000000000000ad2a000000000400a8970100000000000000000000000000bb2a00000100010000030100000000002300000000000000c42a000000000400b6970100000000000000000000000000d12a00000100010000040100000000001000000000000000fc2a000000000400d09701000000000000000000000000000a2b00000100010048040100000000001000000000000000352b0000020004002c980100000000000a000000000000006b2b000000000400e29701000000000000000000000000000000000000000400f09701000000000000000000000000000000000000000400f0970100000000000000000000000000792b00000000040008980100000000000000000000000000872b0000000004001698010000000000000000000000000000000000000004002c98010000000000000000000000000000000000000004002c980100000000000000000000000000000000000000040036980100000000000000000000000000000000000000040036980100000000000000000000000000952b00000000040054980100000000000000000000000000a32b0000000004005e980100000000000000000000000000b12b0000000004006c980100000000000000000000000000000000000000040082980100000000000000000000000000000000000000040082980100000000000000000000000000bf2b000000000400a2980100000000000000000000000000cd2b000000000400ac980100000000000000000000000000db2b000000000400c2980100000000000000000000000000e92b00000100010058040100000000000d000000000000000000000000000400ce980100000000000000000000000000142c000002000400ce98010000000000f4000000000000000000000000000400ce980100000000000000000000000000532c0000000004009a990100000000000000000000000000612c000000000400ae9901000000000000000000000000006f2c000000000400b89901000000000000000000000000000000000000000400c29901000000000000000000000000000000000000000400c29901000000000000000000000000000000000000000400c49901000000000000000000000000000000000000000400dc9901000000000000000000000000007d2c000000000400e29901000000000000000000000000008b2c000001000600e0c9020000000000a800000000000000b32c000000000400ee990100000000000000000000000000c12c000000000400989b0100000000000000000000000000cf2c000000000400da9b0100000000000000000000000000dd2c0000000004000a9d0100000000000000000000000000eb2c000000000400149d0100000000000000000000000000f92c000000000400229d0100000000000000000000000000072d000000000400369d0100000000000000000000000000152d000000000400409d0100000000000000000000000000232d000000000400549d0100000000000000000000000000312d0000000004005c9d01000000000000000000000000003f2d000001000100e0020100000000002000000000000000692d000000000400669d0100000000000000000000000000772d0000000004006e9d0100000000000000000000000000852d000000000400789d0100000000000000000000000000932d000000000400809d01000000000000000000000000000000000000000400969d01000000000000000000000000000000000000000400969d01000000000000000000000000000000000000000400989d01000000000000000000000000000000000000000400b29d0100000000000000000000000000a12d000000000400b29d0100000000000000000000000000af2d000000000400d09d0100000000000000000000000000bd2d0000000004001c9e0100000000000000000000000000cb2d000000000400c49e0100000000000000000000000000d92d00000000040014a10100000000000000000000000000e72d0000000004001ea10100000000000000000000000000f52d0000000004002ca10100000000000000000000000000032e00000000040040a10100000000000000000000000000112e00000000040058a101000000000000000000000000001f2e00000000040060a101000000000000000000000000002d2e0000000004006aa101000000000000000000000000003b2e00000000040072a10100000000000000000000000000000000000000040088a10100000000000000000000000000000000000000040088a1010000000000000000000000000000000000000004008aa10100000000000000000000000000000000000000040098a10100000000000000000000000000492e0000020004005ea20100000000005200000000000000912e000002000400b0a20100000000003400000000000000eb2e0000000004003ca20100000000000000000000000000f92e0000010001007004010000000000190000000000000000000000000004005ea2010000000000000000000000000000000000000004005ea20100000000000000000000000000000000000000040060a20100000000000000000000000000000000000000040066a201000000000000000000000000000000000000000400b0a201000000000000000000000000000000000000000400b0a201000000000000000000000000000000000000000400b2a201000000000000000000000000000000000000000400b4a20100000000000000000000000000022f000002000400e4a201000000000074000000000000000000000000000400e4a201000000000000000000000000000000000000000400e4a201000000000000000000000000000000000000000400e6a201000000000000000000000000000000000000000400eca201000000000000000000000000004d2f000002000400b2c50100000000006200000000000000000000000000040058a30100000000000000000000000000802f00000200040058a30100000000003600000000000000000000000000040058a3010000000000000000000000000000000000000004005aa3010000000000000000000000000000000000000004005ca3010000000000000000000000000000000000000004008ea3010000000000000000000000000000000000000004008ea30100000000000000000000000000000000000000040090a3010000000000000000000000000000000000000004009ca301000000000000000000000000000000000000000400faa301000000000000000000000000000000000000000400faa3010000000000000000000000000000000000000004001ca4010000000000000000000000000000000000000004001ca4010000000000000000000000000000000000000004001ea40100000000000000000000000000000000000000040024a40100000000000000000000000000000000000000040056a40100000000000000000000000000000000000000040056a40100000000000000000000000000000000000000040058a40100000000000000000000000000000000000000040066a40100000000000000000000000000cd2f00000000040082a40100000000000000000000000000db2f000001000100c2040100000000000b000000000000000730000000000400dea40100000000000000000000000000153000000000040038a50100000000000000000000000000000000000000040052a50100000000000000000000000000000000000000040052a50100000000000000000000000000000000000000040094a50100000000000000000000000000233000000200040094a50100000000005000000000000000000000000000040094a50100000000000000000000000000000000000000040096a501000000000000000000000000000000000000000400a2a501000000000000000000000000000000000000000400e4a501000000000000000000000000000631000002000400e4a501000000000074000000000000000000000000000400e4a501000000000000000000000000000000000000000400e6a501000000000000000000000000000000000000000400eea50100000000000000000000000000da31000002000400e2c40100000000005200000000000000863200000000040044a60100000000000000000000000000943200000100010090040100000000001c00000000000000000000000000040058a60100000000000000000000000000000000000000040058a6010000000000000000000000000000000000000004005aa60100000000000000000000000000000000000000040066a601000000000000000000000000000000000000000400bca601000000000000000000000000009d32000002000400bca601000000000082000000000000000000000000000400bca601000000000000000000000000000000000000000400bea601000000000000000000000000000000000000000400c6a6010000000000000000000000000000000000000004003ea7010000000000000000000000000025330000020004003ea7010000000000960100000000000000000000000004003ea70100000000000000000000000000000000000000040040a70100000000000000000000000000000000000000040054a70100000000000000000000000000af33000000000400aca80100000000000000000000000000bd33000000000400b6a80100000000000000000000000000cb33000000000400c0a801000000000000000000000000000000000000000400d4a801000000000000000000000000000000000000000400d4a80100000000000000000000000000000000000000040046a90100000000000000000000000000d93300000200040046a90100000000009200000000000000000000000000040046a90100000000000000000000000000000000000000040048a9010000000000000000000000000000000000000004004aa9010000000000000000000000000034340000000004004ea901000000000000000000000000004234000000000100600101000000000000000000000000004c340000000004005ca90100000000000000000000000000553400000000040062a9010000000000000000000000000063340000010001009b050100000000000f000000000000008e340000000004006ea90100000000000000000000000000973400000000040074a90100000000000000000000000000a53400000100010090050100000000000b00000000000000d03400000000040080a90100000000000000000000000000d93400000000040084a90100000000000000000000000000e73400000100010060050100000000000f0000000000000012350000000004008ca901000000000000000000000000002035000001000100700501000000000020000000000000004b3500000000040098a9010000000000000000000000000054350000000004009ea901000000000000000000000000006235000000000400aea901000000000000000000000000006b35000000000400b2a9010000000000000000000000000079350000010001001d050100000000000700000000000000a435000000000400baa90100000000000000000000000000b23500000100010028050100000000002000000000000000dd3500000200040030c201000000000098000000000000000000000000000400d8a901000000000000000000000000002336000002000400d8a901000000000002000000000000000000000000000400d8a901000000000000000000000000000000000000000400daa901000000000000000000000000000000000000000400daa90100000000000000000000000000000000000000040010aa0100000000000000000000000000000000000000040010aa0100000000000000000000000000000000000000040014aa0100000000000000000000000000000000000000040038aa0100000000000000000000000000623600000000040032ab01000000000000000000000000007036000001000100fd040100000000000f000000000000000000000000000400d0ab01000000000000000000000000009c36000002000400d0ab0100000000007a000000000000000000000000000400d0ab01000000000000000000000000000000000000000400d2ab01000000000000000000000000000000000000000400d6ab010000000000000000000000000000000000000004004aac010000000000000000000000000000000000000004004aac010000000000000000000000000000000000000004004cac0100000000000000000000000000000000000000040050ac01000000000000000000000000000000000000000400ccac0100000000000000000000000000dd36000002000400ccac01000000000060010000000000000000000000000400ccac01000000000000000000000000000000000000000400d0ac01000000000000000000000000000000000000000400f4ac010000000000000000000000000000000000000004002cae010000000000000000000000000000000000000004002cae0100000000000000000000000000000000000000040030ae0100000000000000000000000000000000000000040060ae0100000000000000000000000000193700000000040052af01000000000000000000000000002737000001000100f1040100000000000c00000000000000533700000000040096af01000000000000000000000000006137000000000400b2af01000000000000000000000000006f370000000004005cb001000000000000000000000000007d370000000004008ab001000000000000000000000000008b37000000000400f0b00100000000000000000000000000993700000000040080b10100000000000000000000000000a737000000000400aab10100000000000000000000000000b53700000000040072b20100000000000000000000000000c337000001000100b6040100000000000c00000000000000ee3700000000040092b20100000000000000000000000000fc37000001000100ac040100000000000a000000000000000000000000000400eeb201000000000000000000000000000000000000000400eeb20100000000000000000000000000000000000000040006b30100000000000000000000000000000000000000040006b30100000000000000000000000000000000000000040008b3010000000000000000000000000000000000000004002ab3010000000000000000000000000027380000020004002ab3010000000000040000000000000000000000000004002ab3010000000000000000000000000000000000000004002ab3010000000000000000000000000000000000000004002ab3010000000000000000000000000000000000000004002ab3010000000000000000000000000000000000000004002cb3010000000000000000000000000000000000000004002cb3010000000000000000000000000000000000000004002eb3010000000000000000000000000000000000000004002eb3010000000000000000000000000000000000000004002eb3010000000000000000000000000062380000020004002eb3010000000000020000000000000000000000000004002eb3010000000000000000000000000000000000000004002eb3010000000000000000000000000000000000000004002eb3010000000000000000000000000000000000000004002eb30100000000000000000000000000000000000000040030b30100000000000000000000000000000000000000040030b30100000000000000000000000000ec3800000000050080c90200000000000000000000000000f63800000200040030b30100000000004201000000000000000000000000040030b30100000000000000000000000000000000000000040030b30100000000000000000000000000000000000000040030b30100000000000000000000000000000000000000040032b30100000000000000000000000000000000000000040034b30100000000000000000000000000000000000000040036b30100000000000000000000000000273900000000040042b3010000000000000000000000000035390000010001003006010000000000c80000000000000000000000000004004eb30100000000000000000000000000000000000000040052b30100000000000000000000000000613900000000040056b30100000000000000000000000000000000000000040076b30100000000000000000000000000000000000000040078b30100000000000000000000000000000000000000040086b301000000000000000000000000000000000000000400a0b301000000000000000000000000000000000000000400a0b301000000000000000000000000000000000000000400a2b301000000000000000000000000000000000000000400a2b301000000000000000000000000000000000000000400a6b301000000000000000000000000000000000000000400a6b301000000000000000000000000000000000000000400aab301000000000000000000000000000000000000000400aab301000000000000000000000000000000000000000400b2b301000000000000000000000000000000000000000400b2b301000000000000000000000000000000000000000400b4b301000000000000000000000000000000000000000400b4b301000000000000000000000000000000000000000400bcb301000000000000000000000000000000000000000400bcb301000000000000000000000000000000000000000400beb301000000000000000000000000000000000000000400beb301000000000000000000000000000000000000000400c2b301000000000000000000000000000000000000000400c2b301000000000000000000000000000000000000000400cab301000000000000000000000000000000000000000400cab301000000000000000000000000000000000000000400d0b301000000000000000000000000000000000000000400d4b301000000000000000000000000000000000000000400d8b301000000000000000000000000000000000000000400f4b301000000000000000000000000000000000000000400f8b301000000000000000000000000000000000000000400fab301000000000000000000000000000000000000000400fab301000000000000000000000000000000000000000400fcb301000000000000000000000000000000000000000400fcb30100000000000000000000000000000000000000040008b40100000000000000000000000000000000000000040008b4010000000000000000000000000000000000000004000ab4010000000000000000000000000000000000000004000ab40100000000000000000000000000000000000000040014b40100000000000000000000000000000000000000040014b40100000000000000000000000000000000000000040016b4010000000000000000000000000000000000000004001ab40100000000000000000000000000000000000000040022b40100000000000000000000000000000000000000040022b40100000000000000000000000000000000000000040024b40100000000000000000000000000000000000000040024b4010000000000000000000000000000000000000004002eb40100000000000000000000000000000000000000040030b40100000000000000000000000000000000000000040034b40100000000000000000000000000000000000000040034b40100000000000000000000000000000000000000040036b40100000000000000000000000000000000000000040036b40100000000000000000000000000000000000000040042b40100000000000000000000000000000000000000040042b40100000000000000000000000000000000000000040044b40100000000000000000000000000000000000000040044b4010000000000000000000000000000000000000004004cb4010000000000000000000000000000000000000004004cb40100000000000000000000000000000000000000040050b40100000000000000000000000000000000000000040050b40100000000000000000000000000000000000000040056b40100000000000000000000000000000000000000040056b401000000000000000000000000006f3900000000040058b401000000000000000000000000007d39000001000100300a0100000000000000000000000000000000000000040058b40100000000000000000000000000a83900000200040072b4010000000000e40100000000000000000000000004006cb4010000000000000000000000000000000000000004006eb40100000000000000000000000000000000000000040072b40100000000000000000000000000000000000000040072b40100000000000000000000000000000000000000040072b40100000000000000000000000000000000000000040072b40100000000000000000000000000000000000000040072b40100000000000000000000000000000000000000040074b4010000000000000000000000000000000000000004008eb40100000000000000000000000000000000000000040090b40100000000000000000000000000000000000000040090b4010000000000000000000000000000000000000004009cb4010000000000000000000000000000000000000004009cb401000000000000000000000000000000000000000400a8b401000000000000000000000000000000000000000400acb401000000000000000000000000000000000000000400acb401000000000000000000000000000000000000000400b0b401000000000000000000000000000000000000000400b0b401000000000000000000000000000000000000000400b2b401000000000000000000000000000000000000000400b4b401000000000000000000000000000000000000000400b6b401000000000000000000000000000000000000000400b8b401000000000000000000000000000000000000000400bcb401000000000000000000000000000000000000000400beb401000000000000000000000000000000000000000400beb401000000000000000000000000000000000000000400c2b401000000000000000000000000000000000000000400c2b401000000000000000000000000000000000000000400c6b401000000000000000000000000000000000000000400cab401000000000000000000000000000000000000000400cab401000000000000000000000000000000000000000400ccb401000000000000000000000000000000000000000400ccb401000000000000000000000000000000000000000400d4b401000000000000000000000000000000000000000400d4b401000000000000000000000000000000000000000400d6b401000000000000000000000000000000000000000400d6b401000000000000000000000000000000000000000400d8b401000000000000000000000000000000000000000400d8b401000000000000000000000000000000000000000400dab401000000000000000000000000000000000000000400dab401000000000000000000000000000000000000000400dcb401000000000000000000000000000000000000000400deb401000000000000000000000000000000000000000400e0b401000000000000000000000000000000000000000400e4b401000000000000000000000000000000000000000400e8b401000000000000000000000000000000000000000400e8b401000000000000000000000000000000000000000400eab401000000000000000000000000000000000000000400eab401000000000000000000000000000000000000000400ecb401000000000000000000000000000000000000000400ecb401000000000000000000000000000000000000000400f2b401000000000000000000000000000000000000000400f2b401000000000000000000000000000000000000000400f6b401000000000000000000000000000000000000000400f6b401000000000000000000000000000000000000000400fcb401000000000000000000000000000000000000000400fcb40100000000000000000000000000e13900000200040056b6010000000000560000000000000000000000000004001cb50100000000000000000000000000000000000000040038b5010000000000000000000000000000000000000004003cb50100000000000000000000000000000000000000040062b50100000000000000000000000000000000000000040062b50100000000000000000000000000000000000000040068b50100000000000000000000000000000000000000040068b5010000000000000000000000000000000000000004006cb5010000000000000000000000000000000000000004006cb50100000000000000000000000000000000000000040076b50100000000000000000000000000000000000000040076b5010000000000000000000000000000000000000004007ab5010000000000000000000000000000000000000004007ab5010000000000000000000000000000000000000004007eb5010000000000000000000000000000000000000004007eb50100000000000000000000000000000000000000040092b50100000000000000000000000000000000000000040094b50100000000000000000000000000000000000000040094b5010000000000000000000000000000000000000004009ab5010000000000000000000000000000000000000004009ab5010000000000000000000000000000000000000004009eb5010000000000000000000000000000000000000004009eb501000000000000000000000000000000000000000400aeb501000000000000000000000000000000000000000400aeb501000000000000000000000000000000000000000400b0b501000000000000000000000000000000000000000400b0b501000000000000000000000000000000000000000400b4b501000000000000000000000000000000000000000400b8b501000000000000000000000000000000000000000400bab501000000000000000000000000000000000000000400c0b501000000000000000000000000000000000000000400ccb501000000000000000000000000000000000000000400d0b501000000000000000000000000000000000000000400d0b501000000000000000000000000000000000000000400d2b501000000000000000000000000000000000000000400d2b501000000000000000000000000000000000000000400d4b501000000000000000000000000000000000000000400d4b501000000000000000000000000000000000000000400e0b501000000000000000000000000000000000000000400e0b501000000000000000000000000000000000000000400eab501000000000000000000000000000000000000000400eeb50100000000000000000000000000000000000000040002b60100000000000000000000000000000000000000040010b60100000000000000000000000000000000000000040010b60100000000000000000000000000000000000000040018b60100000000000000000000000000000000000000040018b60100000000000000000000000000000000000000040020b60100000000000000000000000000000000000000040020b60100000000000000000000000000000000000000040030b60100000000000000000000000000000000000000040030b60100000000000000000000000000000000000000040040b60100000000000000000000000000000000000000040042b60100000000000000000000000000000000000000040046b6010000000000000000000000000000000000000004004eb60100000000000000000000000000000000000000040050b60100000000000000000000000000000000000000040050b60100000000000000000000000000000000000000040056b60100000000000000000000000000000000000000040056b60100000000000000000000000000000000000000040056b60100000000000000000000000000000000000000040056b60100000000000000000000000000000000000000040056b60100000000000000000000000000000000000000040056b60100000000000000000000000000000000000000040058b60100000000000000000000000000000000000000040062b60100000000000000000000000000000000000000040072b60100000000000000000000000000000000000000040076b60100000000000000000000000000000000000000040084b60100000000000000000000000000000000000000040086b60100000000000000000000000000000000000000040098b6010000000000000000000000000000000000000004009cb6010000000000000000000000000000000000000004009eb601000000000000000000000000000000000000000400a8b601000000000000000000000000000000000000000400acb601000000000000000000000000000000000000000400acb60100000000000000000000000000283a00000000050088c90200000000000000000000000000323a00000000050090c902000000000000000000000000003c3a000002000400acb601000000000078030000000000000000000000000400acb601000000000000000000000000000000000000000400acb601000000000000000000000000000000000000000400acb601000000000000000000000000000000000000000400aeb601000000000000000000000000000000000000000400aeb601000000000000000000000000000000000000000400aeb601000000000000000000000000000000000000000400c0b601000000000000000000000000000000000000000400c4b601000000000000000000000000000000000000000400c4b601000000000000000000000000000000000000000400c6b601000000000000000000000000000000000000000400c6b601000000000000000000000000000000000000000400ceb601000000000000000000000000000000000000000400ceb601000000000000000000000000000000000000000400d2b601000000000000000000000000000000000000000400d6b601000000000000000000000000000000000000000400dab601000000000000000000000000000000000000000400dab601000000000000000000000000000000000000000400deb601000000000000000000000000000000000000000400deb601000000000000000000000000000000000000000400f0b601000000000000000000000000000000000000000400f0b601000000000000000000000000000000000000000400f4b601000000000000000000000000000000000000000400f4b601000000000000000000000000000000000000000400f6b601000000000000000000000000000000000000000400fab601000000000000000000000000000000000000000400fab601000000000000000000000000000000000000000400feb601000000000000000000000000000000000000000400feb60100000000000000000000000000000000000000040000b70100000000000000000000000000000000000000040000b70100000000000000000000000000000000000000040002b70100000000000000000000000000000000000000040002b70100000000000000000000000000000000000000040006b70100000000000000000000000000000000000000040006b7010000000000000000000000000000000000000004000eb70100000000000000000000000000000000000000040012b70100000000000000000000000000000000000000040016b70100000000000000000000000000000000000000040016b7010000000000000000000000000000000000000004001ab7010000000000000000000000000000000000000004001ab7010000000000000000000000000000000000000004001eb7010000000000000000000000000000000000000004001eb70100000000000000000000000000000000000000040022b70100000000000000000000000000000000000000040026b70100000000000000000000000000000000000000040026b70100000000000000000000000000000000000000040028b7010000000000000000000000000000000000000004002cb70100000000000000000000000000000000000000040030b70100000000000000000000000000000000000000040030b70100000000000000000000000000000000000000040034b70100000000000000000000000000000000000000040038b7010000000000000000000000000000000000000004003cb7010000000000000000000000000000000000000004003cb7010000000000000000000000000000000000000004003eb70100000000000000000000000000000000000000040042b70100000000000000000000000000000000000000040046b70100000000000000000000000000000000000000040046b70100000000000000000000000000000000000000040048b70100000000000000000000000000000000000000040048b7010000000000000000000000000000000000000004004cb7010000000000000000000000000000000000000004004cb7010000000000000000000000000000000000000004006ab7010000000000000000000000000000000000000004006ab7010000000000000000000000000000000000000004006eb7010000000000000000000000000000000000000004006eb70100000000000000000000000000000000000000040072b70100000000000000000000000000000000000000040076b7010000000000000000000000000000000000000004007eb70100000000000000000000000000000000000000040082b70100000000000000000000000000000000000000040086b7010000000000000000000000000000000000000004008ab7010000000000000000000000000000000000000004008eb70100000000000000000000000000000000000000040092b70100000000000000000000000000000000000000040092b70100000000000000000000000000000000000000040096b70100000000000000000000000000000000000000040096b7010000000000000000000000000000000000000004009ab7010000000000000000000000000000000000000004009ab7010000000000000000000000000000000000000004009eb701000000000000000000000000000000000000000400a2b701000000000000000000000000000000000000000400a2b701000000000000000000000000000000000000000400a8b701000000000000000000000000000000000000000400acb701000000000000000000000000000000000000000400aeb701000000000000000000000000000000000000000400aeb701000000000000000000000000000000000000000400b4b701000000000000000000000000000000000000000400b4b701000000000000000000000000000000000000000400b8b701000000000000000000000000000000000000000400b8b701000000000000000000000000000000000000000400bab701000000000000000000000000000000000000000400beb701000000000000000000000000000000000000000400beb701000000000000000000000000000000000000000400c2b701000000000000000000000000000000000000000400c2b701000000000000000000000000000000000000000400cab701000000000000000000000000000000000000000400cab701000000000000000000000000000000000000000400ceb701000000000000000000000000000000000000000400ceb701000000000000000000000000000000000000000400d0b701000000000000000000000000000000000000000400d0b701000000000000000000000000000000000000000400d4b701000000000000000000000000000000000000000400d4b701000000000000000000000000000000000000000400d8b701000000000000000000000000000000000000000400d8b701000000000000000000000000000000000000000400dab701000000000000000000000000000000000000000400dab701000000000000000000000000000000000000000400dcb701000000000000000000000000000000000000000400dcb701000000000000000000000000000000000000000400e0b701000000000000000000000000000000000000000400e4b701000000000000000000000000000000000000000400ecb701000000000000000000000000000000000000000400ecb701000000000000000000000000000000000000000400f0b701000000000000000000000000000000000000000400f2b701000000000000000000000000000000000000000400f2b701000000000000000000000000000000000000000400f6b701000000000000000000000000000000000000000400f6b701000000000000000000000000000000000000000400fab701000000000000000000000000000000000000000400feb701000000000000000000000000000000000000000400feb70100000000000000000000000000000000000000040000b80100000000000000000000000000000000000000040000b80100000000000000000000000000000000000000040008b80100000000000000000000000000000000000000040008b8010000000000000000000000000000000000000004000ab8010000000000000000000000000000000000000004000ab8010000000000000000000000000000000000000004000cb8010000000000000000000000000000000000000004000cb80100000000000000000000000000000000000000040010b80100000000000000000000000000000000000000040010b80100000000000000000000000000000000000000040016b80100000000000000000000000000000000000000040016b8010000000000000000000000000000000000000004001eb8010000000000000000000000000000000000000004001eb80100000000000000000000000000000000000000040024b80100000000000000000000000000000000000000040024b80100000000000000000000000000000000000000040028b80100000000000000000000000000000000000000040028b8010000000000000000000000000000000000000004002ab8010000000000000000000000000000000000000004002eb8010000000000000000000000000000000000000004002eb80100000000000000000000000000000000000000040030b80100000000000000000000000000000000000000040030b80100000000000000000000000000000000000000040038b80100000000000000000000000000000000000000040038b8010000000000000000000000000000000000000004003ab8010000000000000000000000000000000000000004003ab8010000000000000000000000000000000000000004003cb8010000000000000000000000000000000000000004003cb8010000000000000000000000000000000000000004003eb8010000000000000000000000000000000000000004003eb80100000000000000000000000000000000000000040040b80100000000000000000000000000000000000000040040b80100000000000000000000000000000000000000040042b80100000000000000000000000000000000000000040042b80100000000000000000000000000000000000000040048b8010000000000000000000000000000000000000004004cb8010000000000000000000000000000000000000004004cb8010000000000000000000000000000000000000004004eb8010000000000000000000000000000000000000004004eb80100000000000000000000000000000000000000040056b80100000000000000000000000000000000000000040056b80100000000000000000000000000000000000000040058b80100000000000000000000000000000000000000040058b8010000000000000000000000000000000000000004005ab8010000000000000000000000000000000000000004005ab8010000000000000000000000000000000000000004005cb8010000000000000000000000000000000000000004005cb801000000000000000000000000006b3a00000000040060b80100000000000000000000000000793a00000000040068b8010000000000000000000000000000000000000004007eb80100000000000000000000000000000000000000040084b80100000000000000000000000000000000000000040092b80100000000000000000000000000000000000000040092b80100000000000000000000000000000000000000040096b80100000000000000000000000000000000000000040098b8010000000000000000000000000000000000000004009cb8010000000000000000000000000000000000000004009eb8010000000000000000000000000000000000000004009eb801000000000000000000000000000000000000000400a2b801000000000000000000000000000000000000000400a2b801000000000000000000000000000000000000000400a4b801000000000000000000000000000000000000000400a4b801000000000000000000000000000000000000000400a6b801000000000000000000000000000000000000000400a8b801000000000000000000000000000000000000000400a8b801000000000000000000000000000000000000000400aab801000000000000000000000000000000000000000400b4b801000000000000000000000000000000000000000400b8b801000000000000000000000000000000000000000400bcb801000000000000000000000000000000000000000400bcb801000000000000000000000000000000000000000400c0b801000000000000000000000000000000000000000400c0b801000000000000000000000000000000000000000400c6b801000000000000000000000000000000000000000400c6b801000000000000000000000000000000000000000400c8b801000000000000000000000000000000000000000400c8b801000000000000000000000000000000000000000400ccb801000000000000000000000000000000000000000400ceb801000000000000000000000000000000000000000400d0b801000000000000000000000000000000000000000400d0b801000000000000000000000000000000000000000400d4b801000000000000000000000000000000000000000400d6b801000000000000000000000000000000000000000400d8b801000000000000000000000000000000000000000400d8b801000000000000000000000000000000000000000400dab801000000000000000000000000000000000000000400dab801000000000000000000000000000000000000000400deb801000000000000000000000000000000000000000400deb801000000000000000000000000000000000000000400e0b801000000000000000000000000000000000000000400e0b801000000000000000000000000000000000000000400e4b801000000000000000000000000000000000000000400e6b801000000000000000000000000000000000000000400e6b801000000000000000000000000000000000000000400e8b801000000000000000000000000000000000000000400e8b801000000000000000000000000000000000000000400eab801000000000000000000000000000000000000000400eeb801000000000000000000000000000000000000000400f2b801000000000000000000000000000000000000000400f4b801000000000000000000000000000000000000000400f6b801000000000000000000000000000000000000000400f8b801000000000000000000000000000000000000000400f8b801000000000000000000000000000000000000000400fab801000000000000000000000000000000000000000400fab801000000000000000000000000000000000000000400fcb801000000000000000000000000000000000000000400fcb80100000000000000000000000000000000000000040000b90100000000000000000000000000000000000000040000b90100000000000000000000000000000000000000040004b90100000000000000000000000000000000000000040006b90100000000000000000000000000000000000000040008b9010000000000000000000000000000000000000004000cb9010000000000000000000000000000000000000004000cb90100000000000000000000000000000000000000040010b90100000000000000000000000000000000000000040010b90100000000000000000000000000000000000000040012b90100000000000000000000000000000000000000040012b90100000000000000000000000000000000000000040018b90100000000000000000000000000000000000000040018b9010000000000000000000000000000000000000004001cb90100000000000000000000000000000000000000040020b90100000000000000000000000000000000000000040024b9010000000000000000000000000000000000000004002ab90100000000000000000000000000000000000000040030b90100000000000000000000000000000000000000040030b90100000000000000000000000000000000000000040032b90100000000000000000000000000000000000000040032b90100000000000000000000000000000000000000040034b90100000000000000000000000000000000000000040034b90100000000000000000000000000000000000000040038b9010000000000000000000000000000000000000004003ab9010000000000000000000000000000000000000004003cb90100000000000000000000000000000000000000040040b90100000000000000000000000000000000000000040040b90100000000000000000000000000000000000000040042b90100000000000000000000000000000000000000040042b90100000000000000000000000000000000000000040044b90100000000000000000000000000000000000000040044b90100000000000000000000000000000000000000040048b90100000000000000000000000000000000000000040048b9010000000000000000000000000000000000000004004ab9010000000000000000000000000000000000000004004ab9010000000000000000000000000000000000000004004eb90100000000000000000000000000000000000000040050b90100000000000000000000000000000000000000040054b90100000000000000000000000000000000000000040056b90100000000000000000000000000000000000000040056b9010000000000000000000000000000000000000004005ab9010000000000000000000000000000000000000004005ab9010000000000000000000000000000000000000004005cb9010000000000000000000000000000000000000004005cb9010000000000000000000000000000000000000004005eb9010000000000000000000000000000000000000004005eb90100000000000000000000000000000000000000040062b90100000000000000000000000000000000000000040062b90100000000000000000000000000000000000000040068b90100000000000000000000000000000000000000040068b9010000000000000000000000000000000000000004006cb9010000000000000000000000000000000000000004006cb90100000000000000000000000000000000000000040072b90100000000000000000000000000000000000000040072b90100000000000000000000000000000000000000040098b90100000000000000000000000000000000000000040098b9010000000000000000000000000000000000000004009cb901000000000000000000000000000000000000000400a0b901000000000000000000000000000000000000000400a2b901000000000000000000000000000000000000000400a8b901000000000000000000000000000000000000000400b6b901000000000000000000000000000000000000000400bab901000000000000000000000000000000000000000400bab901000000000000000000000000000000000000000400bcb901000000000000000000000000000000000000000400bcb901000000000000000000000000000000000000000400beb901000000000000000000000000000000000000000400beb901000000000000000000000000000000000000000400cab901000000000000000000000000000000000000000400cab901000000000000000000000000000000000000000400d4b901000000000000000000000000000000000000000400d8b901000000000000000000000000000000000000000400e6b901000000000000000000000000000000000000000400e6b901000000000000000000000000000000000000000400eeb901000000000000000000000000000000000000000400eeb901000000000000000000000000000000000000000400f2b901000000000000000000000000000000000000000400f2b901000000000000000000000000000000000000000400f6b901000000000000000000000000000000000000000400f6b90100000000000000000000000000000000000000040006ba0100000000000000000000000000000000000000040008ba0100000000000000000000000000000000000000040008ba010000000000000000000000000000000000000004000cba010000000000000000000000000000000000000004000cba0100000000000000000000000000000000000000040020ba0100000000000000000000000000000000000000040024ba0100000000000000000000000000000000000000040024ba0100000000000000000000000000000000000000040024ba0100000000000000000000000000000000000000040024ba0100000000000000000000000000000000000000040024ba0100000000000000000000000000000000000000040026ba0100000000000000000000000000000000000000040026ba0100000000000000000000000000000000000000040028ba0100000000000000000000000000000000000000040032ba0100000000000000000000000000000000000000040032ba0100000000000000000000000000873a00000200040032ba0100000000007e01000000000000000000000000040032ba0100000000000000000000000000000000000000040032ba0100000000000000000000000000000000000000040032ba0100000000000000000000000000000000000000040034ba0100000000000000000000000000000000000000040044ba010000000000000000000000000000000000000004004aba010000000000000000000000000000000000000004004aba0100000000000000000000000000000000000000040052ba0100000000000000000000000000000000000000040052ba0100000000000000000000000000000000000000040056ba0100000000000000000000000000000000000000040056ba010000000000000000000000000000000000000004005eba010000000000000000000000000000000000000004005eba0100000000000000000000000000000000000000040060ba0100000000000000000000000000000000000000040064ba0100000000000000000000000000000000000000040064ba0100000000000000000000000000000000000000040068ba010000000000000000000000000000000000000004006cba0100000000000000000000000000ae3a00000000040086ba010000000000000000000000000000000000000004008eba010000000000000000000000000000000000000004008eba0100000000000000000000000000000000000000040090ba0100000000000000000000000000000000000000040092ba0100000000000000000000000000000000000000040096ba010000000000000000000000000000000000000004009aba01000000000000000000000000000000000000000400a0ba01000000000000000000000000000000000000000400a0ba01000000000000000000000000000000000000000400a2ba01000000000000000000000000000000000000000400a4ba01000000000000000000000000000000000000000400a8ba01000000000000000000000000000000000000000400acba01000000000000000000000000000000000000000400aeba01000000000000000000000000000000000000000400aeba01000000000000000000000000000000000000000400b2ba01000000000000000000000000000000000000000400b2ba01000000000000000000000000000000000000000400b4ba01000000000000000000000000000000000000000400baba01000000000000000000000000000000000000000400baba01000000000000000000000000000000000000000400c0ba01000000000000000000000000000000000000000400c0ba01000000000000000000000000000000000000000400caba01000000000000000000000000000000000000000400ceba01000000000000000000000000000000000000000400d0ba01000000000000000000000000000000000000000400d2ba01000000000000000000000000000000000000000400d2ba01000000000000000000000000000000000000000400d4ba01000000000000000000000000000000000000000400d8ba01000000000000000000000000000000000000000400e0ba01000000000000000000000000000000000000000400e0ba01000000000000000000000000000000000000000400e6ba01000000000000000000000000000000000000000400e6ba01000000000000000000000000000000000000000400f0ba01000000000000000000000000000000000000000400f4ba01000000000000000000000000000000000000000400f6ba01000000000000000000000000000000000000000400f8ba01000000000000000000000000000000000000000400f8ba01000000000000000000000000000000000000000400faba01000000000000000000000000000000000000000400feba0100000000000000000000000000000000000000040000bb0100000000000000000000000000000000000000040000bb0100000000000000000000000000000000000000040004bb0100000000000000000000000000000000000000040004bb0100000000000000000000000000000000000000040006bb0100000000000000000000000000000000000000040008bb010000000000000000000000000000000000000004000cbb010000000000000000000000000000000000000004000cbb010000000000000000000000000000000000000004000ebb010000000000000000000000000000000000000004000ebb010000000000000000000000000000000000000004001ebb010000000000000000000000000000000000000004001ebb0100000000000000000000000000000000000000040022bb0100000000000000000000000000000000000000040022bb0100000000000000000000000000000000000000040026bb010000000000000000000000000000000000000004002ebb0100000000000000000000000000000000000000040040bb0100000000000000000000000000000000000000040040bb0100000000000000000000000000000000000000040042bb0100000000000000000000000000000000000000040044bb0100000000000000000000000000000000000000040048bb010000000000000000000000000000000000000004004cbb0100000000000000000000000000000000000000040052bb0100000000000000000000000000000000000000040052bb0100000000000000000000000000000000000000040054bb0100000000000000000000000000000000000000040058bb010000000000000000000000000000000000000004005cbb010000000000000000000000000000000000000004005cbb010000000000000000000000000000000000000004005ebb010000000000000000000000000000000000000004005ebb0100000000000000000000000000000000000000040068bb0100000000000000000000000000000000000000040068bb010000000000000000000000000000000000000004006cbb010000000000000000000000000000000000000004006cbb0100000000000000000000000000000000000000040072bb0100000000000000000000000000000000000000040072bb0100000000000000000000000000000000000000040074bb0100000000000000000000000000000000000000040078bb0100000000000000000000000000000000000000040078bb010000000000000000000000000000000000000004007cbb010000000000000000000000000000000000000004007cbb0100000000000000000000000000000000000000040080bb0100000000000000000000000000000000000000040080bb0100000000000000000000000000000000000000040084bb0100000000000000000000000000000000000000040084bb0100000000000000000000000000000000000000040088bb0100000000000000000000000000000000000000040090bb0100000000000000000000000000000000000000040096bb010000000000000000000000000000000000000004009cbb01000000000000000000000000000000000000000400acbb01000000000000000000000000000000000000000400b0bb01000000000000000000000000000000000000000400b0bb0100000000000000000000000000bc3a000002000400b0bb01000000000012000000000000000000000000000400b0bb01000000000000000000000000000000000000000400b0bb01000000000000000000000000000000000000000400b0bb01000000000000000000000000000000000000000400b0bb0100000000000000000000000000163b000000000400b6bb0100000000000000000000000000243b000001000100cd050100000000000b000000000000000000000000000400c2bb01000000000000000000000000000000000000000400c2bb01000000000000000000000000000000000000000400c2bb0100000000000000000000000000503b000002000400c2bb01000000000012000000000000000000000000000400c2bb01000000000000000000000000000000000000000400c2bb01000000000000000000000000000000000000000400c2bb01000000000000000000000000000000000000000400c2bb0100000000000000000000000000ad3b000000000400c8bb0100000000000000000000000000bb3b000001000100d8050100000000000e000000000000000000000000000400d4bb01000000000000000000000000000000000000000400d4bb01000000000000000000000000000000000000000400d4bb01000000000000000000000000000000000000000400d4bb01000000000000000000000000000000000000000400d4bb01000000000000000000000000000000000000000400d4bb01000000000000000000000000000000000000000400d6bb01000000000000000000000000000000000000000400d6bb01000000000000000000000000000000000000000400d8bb01000000000000000000000000000000000000000400e2bb01000000000000000000000000000000000000000400e2bb01000000000000000000000000000000000000000400e2bb01000000000000000000000000000000000000000400e2bb01000000000000000000000000000000000000000400e2bb01000000000000000000000000000000000000000400e4bb01000000000000000000000000000000000000000400e4bb01000000000000000000000000000000000000000400e4bb01000000000000000000000000000000000000000400e6bb01000000000000000000000000000000000000000400f0bb01000000000000000000000000000000000000000400f0bb01000000000000000000000000000000000000000400f0bb01000000000000000000000000000000000000000400f0bb01000000000000000000000000000000000000000400f0bb01000000000000000000000000000000000000000400f0bb01000000000000000000000000000000000000000400f2bb01000000000000000000000000000000000000000400f2bb01000000000000000000000000000000000000000400f4bb01000000000000000000000000000000000000000400febb01000000000000000000000000000000000000000400febb0100000000000000000000000000e73b000002000400febb01000000000070000000000000000000000000000400febb01000000000000000000000000000000000000000400febb01000000000000000000000000000000000000000400febb0100000000000000000000000000000000000000040000bc0100000000000000000000000000000000000000040002bc0100000000000000000000000000000000000000040004bc0100000000000000000000000000000000000000040004bc010000000000000000000000000000000000000004000cbc010000000000000000000000000000000000000004000cbc0100000000000000000000000000000000000000040014bc0100000000000000000000000000000000000000040014bc0100000000000000000000000000000000000000040016bc0100000000000000000000000000000000000000040016bc010000000000000000000000000000000000000004001abc010000000000000000000000000000000000000004001abc0100000000000000000000000000000000000000040022bc0100000000000000000000000000000000000000040024bc0100000000000000000000000000000000000000040024bc010000000000000000000000000000000000000004002cbc010000000000000000000000000000000000000004002cbc0100000000000000000000000000000000000000040030bc0100000000000000000000000000000000000000040030bc010000000000000000000000000000000000000004003abc010000000000000000000000000000000000000004003abc0100000000000000000000000000000000000000040044bc0100000000000000000000000000473c00000000040044bc0100000000000000000000000000553c0000010001002e060100000000000200000000000000000000000000040044bc010000000000000000000000000000000000000004005abc010000000000000000000000000000000000000004005abc010000000000000000000000000000000000000004005cbc0100000000000000000000000000000000000000040060bc0100000000000000000000000000000000000000040060bc010000000000000000000000000000000000000004006ebc010000000000000000000000000000000000000004006ebc010000000000000000000000000000000000000004006ebc0100000000000000000000000000813c00000000050098c902000000000000000000000000008c3c000000000500a0c90200000000000000000000000000973c000000000500a8c90200000000000000000000000000a23c0000020004006ebc010000000000bc0100000000000000000000000004006ebc010000000000000000000000000000000000000004006ebc010000000000000000000000000000000000000004006ebc0100000000000000000000000000000000000000040070bc010000000000000000000000000000000000000004008abc01000000000000000000000000000a3d00000000040094bc0100000000000000000000000000183d0000000004009cbc0100000000000000000000000000263d000000000400a4bc01000000000000000000000000000000000000000400b4bc01000000000000000000000000000000000000000400b4bc0100000000000000000000000000343d000000000400bcbc01000000000000000000000000000000000000000400ccbc01000000000000000000000000000000000000000400ccbc01000000000000000000000000000000000000000400d0bc01000000000000000000000000000000000000000400d0bc01000000000000000000000000000000000000000400dabc01000000000000000000000000000000000000000400dabc01000000000000000000000000000000000000000400debc01000000000000000000000000000000000000000400ecbc01000000000000000000000000000000000000000400ecbc01000000000000000000000000000000000000000400f4bc01000000000000000000000000000000000000000400f4bc01000000000000000000000000000000000000000400febc01000000000000000000000000000000000000000400febc0100000000000000000000000000000000000000040006bd0100000000000000000000000000000000000000040006bd010000000000000000000000000000000000000004000cbd010000000000000000000000000000000000000004000cbd0100000000000000000000000000000000000000040010bd0100000000000000000000000000000000000000040012bd010000000000000000000000000000000000000004001ebd0100000000000000000000000000000000000000040020bd0100000000000000000000000000000000000000040026bd0100000000000000000000000000000000000000040026bd010000000000000000000000000000000000000004002ebd0100000000000000000000000000000000000000040032bd0100000000000000000000000000000000000000040032bd0100000000000000000000000000000000000000040040bd0100000000000000000000000000000000000000040046bd010000000000000000000000000000000000000004004abd010000000000000000000000000000000000000004004abd010000000000000000000000000000000000000004004ebd010000000000000000000000000000000000000004004ebd0100000000000000000000000000000000000000040054bd0100000000000000000000000000000000000000040056bd0100000000000000000000000000000000000000040056bd0100000000000000000000000000000000000000040058bd0100000000000000000000000000000000000000040058bd0100000000000000000000000000000000000000040060bd0100000000000000000000000000000000000000040060bd010000000000000000000000000000000000000004006abd010000000000000000000000000000000000000004006cbd010000000000000000000000000000000000000004006cbd010000000000000000000000000000000000000004006ebd010000000000000000000000000000000000000004006ebd0100000000000000000000000000000000000000040076bd0100000000000000000000000000000000000000040076bd0100000000000000000000000000000000000000040078bd010000000000000000000000000000000000000004007ebd010000000000000000000000000000000000000004007ebd010000000000000000000000000000000000000004008abd010000000000000000000000000000000000000004008cbd0100000000000000000000000000000000000000040090bd0100000000000000000000000000000000000000040090bd0100000000000000000000000000000000000000040094bd0100000000000000000000000000000000000000040098bd010000000000000000000000000000000000000004009ebd010000000000000000000000000000000000000004009ebd01000000000000000000000000000000000000000400aabd01000000000000000000000000000000000000000400b2bd01000000000000000000000000000000000000000400b2bd01000000000000000000000000000000000000000400b4bd01000000000000000000000000000000000000000400b6bd01000000000000000000000000000000000000000400bebd01000000000000000000000000000000000000000400bebd01000000000000000000000000000000000000000400c0bd01000000000000000000000000000000000000000400c0bd01000000000000000000000000000000000000000400c4bd01000000000000000000000000000000000000000400c4bd01000000000000000000000000000000000000000400c8bd01000000000000000000000000000000000000000400c8bd01000000000000000000000000000000000000000400dcbd01000000000000000000000000000000000000000400e2bd01000000000000000000000000000000000000000400f0bd01000000000000000000000000000000000000000400f8bd01000000000000000000000000000000000000000400f8bd01000000000000000000000000000000000000000400fcbd01000000000000000000000000000000000000000400fcbd010000000000000000000000000000000000000004000cbe0100000000000000000000000000000000000000040026be010000000000000000000000000000000000000004002abe010000000000000000000000000000000000000004002abe0100000000000000000000000000423d0000020004002abe010000000000b40000000000000000000000000004002abe010000000000000000000000000000000000000004002abe010000000000000000000000000000000000000004002abe010000000000000000000000000000000000000004002cbe010000000000000000000000000000000000000004002ebe0100000000000000000000000000000000000000040036be0100000000000000000000000000000000000000040038be0100000000000000000000000000000000000000040038be010000000000000000000000000000000000000004003cbe010000000000000000000000000000000000000004003cbe0100000000000000000000000000000000000000040044be0100000000000000000000000000000000000000040044be010000000000000000000000000000000000000004004abe010000000000000000000000000000000000000004004abe010000000000000000000000000000000000000004004ebe0100000000000000000000000000000000000000040056be010000000000000000000000000000000000000004005abe0100000000000000000000000000000000000000040066be0100000000000000000000000000000000000000040066be010000000000000000000000000000000000000004006cbe010000000000000000000000000000000000000004006cbe0100000000000000000000000000000000000000040070be0100000000000000000000000000000000000000040078be010000000000000000000000000000000000000004007ebe0100000000000000000000000000000000000000040086be010000000000000000000000000000000000000004008abe0100000000000000000000000000000000000000040096be010000000000000000000000000000000000000004009cbe01000000000000000000000000000000000000000400a4be01000000000000000000000000000000000000000400aabe01000000000000000000000000000000000000000400b2be01000000000000000000000000000000000000000400b8be01000000000000000000000000000000000000000400c0be01000000000000000000000000000000000000000400c4be01000000000000000000000000000000000000000400cebe01000000000000000000000000000000000000000400cebe01000000000000000000000000000000000000000400d8be01000000000000000000000000000000000000000400dabe01000000000000000000000000000000000000000400debe01000000000000000000000000000000000000000400debe0100000000000000000000000000753d000002000400debe01000000000038000000000000000000000000000400debe01000000000000000000000000000000000000000400debe01000000000000000000000000000000000000000400debe01000000000000000000000000000000000000000400e0be01000000000000000000000000000000000000000400e0be01000000000000000000000000000000000000000400e2be0100000000000000000000000000a63d000000000400fcbe0100000000000000000000000000b43d000001000100f8060100000000003000000000000000000000000000040010bf0100000000000000000000000000000000000000040012bf0100000000000000000000000000000000000000040016bf0100000000000000000000000000000000000000040016bf0100000000000000000000000000e03d00000200040016bf0100000000000a00000000000000000000000000040016bf0100000000000000000000000000000000000000040016bf0100000000000000000000000000000000000000040016bf0100000000000000000000000000000000000000040016bf0100000000000000000000000000000000000000040020bf0100000000000000000000000000000000000000040020bf0100000000000000000000000000363e00000200040020bf010000000000b600000000000000000000000000040020bf0100000000000000000000000000000000000000040020bf0100000000000000000000000000000000000000040020bf0100000000000000000000000000000000000000040022bf0100000000000000000000000000000000000000040022bf0100000000000000000000000000000000000000040024bf010000000000000000000000000000000000000004002ebf010000000000000000000000000000000000000004002ebf0100000000000000000000000000000000000000040030bf0100000000000000000000000000000000000000040030bf0100000000000000000000000000000000000000040034bf0100000000000000000000000000000000000000040034bf010000000000000000000000000000000000000004003cbf010000000000000000000000000000000000000004003cbf0100000000000000000000000000000000000000040042bf0100000000000000000000000000000000000000040042bf0100000000000000000000000000000000000000040046bf010000000000000000000000000000000000000004004ebf0100000000000000000000000000000000000000040052bf010000000000000000000000000000000000000004005ebf010000000000000000000000000000000000000004005ebf0100000000000000000000000000000000000000040064bf0100000000000000000000000000000000000000040064bf0100000000000000000000000000000000000000040068bf0100000000000000000000000000000000000000040070bf0100000000000000000000000000000000000000040076bf010000000000000000000000000000000000000004007ebf0100000000000000000000000000000000000000040082bf010000000000000000000000000000000000000004008ebf0100000000000000000000000000000000000000040094bf010000000000000000000000000000000000000004009cbf01000000000000000000000000000000000000000400a2bf01000000000000000000000000000000000000000400aabf01000000000000000000000000000000000000000400b0bf01000000000000000000000000000000000000000400b8bf01000000000000000000000000000000000000000400bcbf01000000000000000000000000000000000000000400c6bf01000000000000000000000000000000000000000400c6bf01000000000000000000000000000000000000000400d0bf01000000000000000000000000000000000000000400d0bf01000000000000000000000000000000000000000400d2bf01000000000000000000000000000000000000000400d6bf01000000000000000000000000000000000000000400d6bf01000000000000000000000000008e3e000002000400d6bf0100000000003a000000000000000000000000000400d6bf01000000000000000000000000000000000000000400d6bf01000000000000000000000000000000000000000400d6bf01000000000000000000000000000000000000000400d8bf01000000000000000000000000000000000000000400d8bf01000000000000000000000000000000000000000400dabf0100000000000000000000000000e43e000000000400f6bf01000000000000000000000000000000000000000400f6bf01000000000000000000000000000000000000000400f6bf010000000000000000000000000000000000000004000ac0010000000000000000000000000000000000000004000ac0010000000000000000000000000000000000000004000cc00100000000000000000000000000000000000000040010c00100000000000000000000000000000000000000040010c00100000000000000000000000000f23e00000200040010c00100000000002001000000000000000000000000040010c00100000000000000000000000000000000000000040010c00100000000000000000000000000000000000000040010c00100000000000000000000000000000000000000040012c00100000000000000000000000000000000000000040020c00100000000000000000000000000000000000000040022c00100000000000000000000000000000000000000040026c00100000000000000000000000000000000000000040026c00100000000000000000000000000000000000000040028c00100000000000000000000000000000000000000040028c00100000000000000000000000000000000000000040030c00100000000000000000000000000000000000000040034c00100000000000000000000000000000000000000040034c00100000000000000000000000000000000000000040038c00100000000000000000000000000000000000000040038c0010000000000000000000000000000000000000004003cc0010000000000000000000000000000000000000004003cc00100000000000000000000000000000000000000040040c00100000000000000000000000000000000000000040040c00100000000000000000000000000000000000000040044c00100000000000000000000000000000000000000040044c00100000000000000000000000000000000000000040046c0010000000000000000000000000000000000000004004ac001000000000000000000000000002e3f0000000004004ec001000000000000000000000000003c3f0000010001002606010000000000020000000000000000000000000004004ec00100000000000000000000000000000000000000040058c0010000000000000000000000000000000000000004005cc0010000000000000000000000000000000000000004005cc00100000000000000000000000000683f00000000040066c00100000000000000000000000000763f00000100010028060100000000000200000000000000000000000000040072c00100000000000000000000000000000000000000040072c00100000000000000000000000000000000000000040074c00100000000000000000000000000a23f0000000004007ac00100000000000000000000000000b03f0000010001002a060100000000000100000000000000000000000000040082c00100000000000000000000000000000000000000040082c0010000000000000000000000000000000000000004008cc0010000000000000000000000000000000000000004008cc0010000000000000000000000000000000000000004008ec0010000000000000000000000000000000000000004008ec00100000000000000000000000000000000000000040092c00100000000000000000000000000000000000000040092c00100000000000000000000000000000000000000040094c00100000000000000000000000000000000000000040094c001000000000000000000000000000000000000000400a0c001000000000000000000000000000000000000000400a0c001000000000000000000000000000000000000000400a4c001000000000000000000000000000000000000000400a4c001000000000000000000000000000000000000000400a6c001000000000000000000000000000000000000000400aac001000000000000000000000000000000000000000400aac001000000000000000000000000000000000000000400b2c001000000000000000000000000000000000000000400b2c001000000000000000000000000000000000000000400bcc001000000000000000000000000000000000000000400bcc001000000000000000000000000000000000000000400c0c001000000000000000000000000000000000000000400c4c001000000000000000000000000000000000000000400ccc001000000000000000000000000000000000000000400d4c001000000000000000000000000000000000000000400e8c001000000000000000000000000000000000000000400e8c001000000000000000000000000000000000000000400ecc00100000000000000000000000000dc3f000000000400ecc00100000000000000000000000000ea3f000001000100e80501000000000030000000000000000000000000000400ecc001000000000000000000000000000000000000000400f6c001000000000000000000000000000000000000000400f6c001000000000000000000000000000000000000000400fec001000000000000000000000000000000000000000400fec00100000000000000000000000000164000000000040004c10100000000000000000000000000244000000100010024060100000000000200000000000000000000000000040010c10100000000000000000000000000000000000000040010c10100000000000000000000000000000000000000040012c10100000000000000000000000000000000000000040012c10100000000000000000000000000000000000000040016c1010000000000000000000000000000000000000004001cc1010000000000000000000000000000000000000004002cc10100000000000000000000000000000000000000040030c10100000000000000000000000000000000000000040030c10100000000000000000000000000504000000200040030c10100000000000001000000000000000000000000040030c10100000000000000000000000000000000000000040030c10100000000000000000000000000000000000000040030c10100000000000000000000000000000000000000040032c10100000000000000000000000000000000000000040040c10100000000000000000000000000000000000000040042c10100000000000000000000000000000000000000040042c1010000000000000000000000000000000000000004004ac1010000000000000000000000000000000000000004004ac1010000000000000000000000000000000000000004004cc1010000000000000000000000000000000000000004004cc10100000000000000000000000000000000000000040050c10100000000000000000000000000000000000000040054c10100000000000000000000000000000000000000040054c10100000000000000000000000000000000000000040064c10100000000000000000000000000000000000000040068c1010000000000000000000000000000000000000004006cc1010000000000000000000000000000000000000004006cc10100000000000000000000000000000000000000040070c10100000000000000000000000000000000000000040070c10100000000000000000000000000000000000000040074c10100000000000000000000000000000000000000040074c10100000000000000000000000000000000000000040078c10100000000000000000000000000000000000000040078c1010000000000000000000000000000000000000004007cc1010000000000000000000000000000000000000004007cc1010000000000000000000000000000000000000004007ec10100000000000000000000000000000000000000040080c10100000000000000000000000000000000000000040080c1010000000000000000000000000089400000000004008ac10100000000000000000000000000000000000000040098c10100000000000000000000000000000000000000040098c1010000000000000000000000000000000000000004009ac101000000000000000000000000000000000000000400a4c101000000000000000000000000000000000000000400a6c101000000000000000000000000000000000000000400a6c101000000000000000000000000009740000000000400b0c10100000000000000000000000000a5400000010001002c0601000000000001000000000000000000000000000400bec101000000000000000000000000000000000000000400bec101000000000000000000000000000000000000000400c0c101000000000000000000000000000000000000000400c0c101000000000000000000000000000000000000000400c4c101000000000000000000000000000000000000000400c4c101000000000000000000000000000000000000000400c6c101000000000000000000000000000000000000000400cac101000000000000000000000000000000000000000400cac101000000000000000000000000000000000000000400d2c101000000000000000000000000000000000000000400d2c101000000000000000000000000000000000000000400dcc101000000000000000000000000000000000000000400dcc101000000000000000000000000000000000000000400e0c101000000000000000000000000000000000000000400e4c101000000000000000000000000000000000000000400ecc101000000000000000000000000000000000000000400f4c10100000000000000000000000000d14000000000040008c20100000000000000000000000000000000000000040012c20100000000000000000000000000000000000000040012c2010000000000000000000000000000000000000004001ac2010000000000000000000000000000000000000004001ac20100000000000000000000000000df4000000000040020c20100000000000000000000000000000000000000040030c20100000000000000000000000000000000000000040030c20100000000000000000000000000000000000000040030c20100000000000000000000000000000000000000040030c20100000000000000000000000000000000000000040030c20100000000000000000000000000000000000000040030c20100000000000000000000000000000000000000040032c2010000000000000000000000000000000000000004003ac2010000000000000000000000000000000000000004003cc2010000000000000000000000000000000000000004003cc20100000000000000000000000000000000000000040048c20100000000000000000000000000000000000000040048c20100000000000000000000000000000000000000040054c20100000000000000000000000000000000000000040054c20100000000000000000000000000000000000000040062c20100000000000000000000000000000000000000040062c20100000000000000000000000000000000000000040064c20100000000000000000000000000000000000000040068c2010000000000000000000000000000000000000004006ac2010000000000000000000000000000000000000004006cc2010000000000000000000000000000000000000004006cc2010000000000000000000000000000000000000004006ec2010000000000000000000000000000000000000004006ec20100000000000000000000000000000000000000040078c2010000000000000000000000000000000000000004007ac20100000000000000000000000000000000000000040082c20100000000000000000000000000000000000000040082c20100000000000000000000000000000000000000040088c20100000000000000000000000000000000000000040088c2010000000000000000000000000000000000000004008ac2010000000000000000000000000000000000000004008ac20100000000000000000000000000ed4000000000040090c20100000000000000000000000000fb400000010001002b06010000000000010000000000000000000000000004009ec2010000000000000000000000000000000000000004009ec201000000000000000000000000000000000000000400a0c201000000000000000000000000000000000000000400a0c201000000000000000000000000002741000000000400a6c201000000000000000000000000003541000001000100cc0501000000000001000000000000000000000000000400b6c201000000000000000000000000000000000000000400b6c201000000000000000000000000000000000000000400bac201000000000000000000000000000000000000000400bac201000000000000000000000000000000000000000400c4c201000000000000000000000000000000000000000400c8c201000000000000000000000000000000000000000400c8c201000000000000000000000000000000000000000400c8c201000000000000000000000000000000000000000400c8c201000000000000000000000000000000000000000400c8c201000000000000000000000000000000000000000400cac201000000000000000000000000000000000000000400cac201000000000000000000000000000000000000000400ccc201000000000000000000000000000000000000000400d6c201000000000000000000000000000000000000000400d6c201000000000000000000000000006141000002000400d6c201000000000072000000000000000000000000000400d6c201000000000000000000000000000000000000000400d6c201000000000000000000000000000000000000000400d6c201000000000000000000000000000000000000000400d8c201000000000000000000000000000000000000000400dac201000000000000000000000000000000000000000400dcc201000000000000000000000000000000000000000400dcc201000000000000000000000000000000000000000400e4c201000000000000000000000000000000000000000400e4c201000000000000000000000000000000000000000400f0c201000000000000000000000000000000000000000400f0c201000000000000000000000000000000000000000400f2c201000000000000000000000000000000000000000400f2c201000000000000000000000000000000000000000400f6c201000000000000000000000000000000000000000400f6c201000000000000000000000000000000000000000400fec201000000000000000000000000000000000000000400fec20100000000000000000000000000000000000000040006c30100000000000000000000000000000000000000040006c3010000000000000000000000000000000000000004000ac3010000000000000000000000000000000000000004000ac30100000000000000000000000000000000000000040014c30100000000000000000000000000000000000000040014c3010000000000000000000000000000000000000004001ec30100000000000000000000000000c0410000000004001ec3010000000000000000000000000000000000000004001ec30100000000000000000000000000000000000000040034c30100000000000000000000000000000000000000040034c30100000000000000000000000000000000000000040036c3010000000000000000000000000000000000000004003ac3010000000000000000000000000000000000000004003ac30100000000000000000000000000000000000000040048c30100000000000000000000000000000000000000040048c30100000000000000000000000000000000000000040048c30100000000000000000000000000ce4100000200040048c30100000000007200000000000000000000000000040048c30100000000000000000000000000000000000000040048c30100000000000000000000000000000000000000040048c3010000000000000000000000000000000000000004004ac3010000000000000000000000000000000000000004004cc3010000000000000000000000000000000000000004004ec3010000000000000000000000000000000000000004004ec30100000000000000000000000000000000000000040056c30100000000000000000000000000000000000000040056c30100000000000000000000000000000000000000040062c30100000000000000000000000000000000000000040062c30100000000000000000000000000000000000000040064c30100000000000000000000000000000000000000040064c30100000000000000000000000000000000000000040068c30100000000000000000000000000000000000000040068c30100000000000000000000000000000000000000040070c30100000000000000000000000000000000000000040070c30100000000000000000000000000000000000000040078c30100000000000000000000000000000000000000040078c3010000000000000000000000000000000000000004007cc3010000000000000000000000000000000000000004007cc30100000000000000000000000000000000000000040086c30100000000000000000000000000000000000000040086c30100000000000000000000000000000000000000040090c301000000000000000000000000002d4200000000040090c30100000000000000000000000000000000000000040090c301000000000000000000000000000000000000000400a6c301000000000000000000000000000000000000000400a6c301000000000000000000000000000000000000000400a8c301000000000000000000000000000000000000000400acc301000000000000000000000000000000000000000400acc301000000000000000000000000000000000000000400bac301000000000000000000000000000000000000000400bac301000000000000000000000000000000000000000400bac301000000000000000000000000003b42000002000400bac301000000000016000000000000000000000000000400bac301000000000000000000000000000000000000000400bac301000000000000000000000000008342000000000400bac301000000000000000000000000000000000000000400bac301000000000000000000000000009142000001000100280701000000000002000000000000000000000000000400bac301000000000000000000000000000000000000000400d0c301000000000000000000000000000000000000000400d0c301000000000000000000000000000000000000000400d0c30100000000000000000000000000bd42000002000400d0c3010000000000a2000000000000000000000000000400d0c301000000000000000000000000000000000000000400d0c301000000000000000000000000000000000000000400d0c301000000000000000000000000000000000000000400d2c301000000000000000000000000000000000000000400d8c301000000000000000000000000000000000000000400dac301000000000000000000000000000000000000000400dac301000000000000000000000000000000000000000400dcc301000000000000000000000000000000000000000400dcc301000000000000000000000000000000000000000400dec301000000000000000000000000000000000000000400dec301000000000000000000000000001e43000000000400e2c301000000000000000000000000002c43000001000100500701000000000011000000000000000000000000000400eec301000000000000000000000000000000000000000400eec301000000000000000000000000000000000000000400fac301000000000000000000000000005843000000000400fac301000000000000000000000000006643000001000100300701000000000020000000000000000000000000000400fac3010000000000000000000000000000000000000004000ec4010000000000000000000000000000000000000004000ec40100000000000000000000000000000000000000040010c40100000000000000000000000000000000000000040014c40100000000000000000000000000000000000000040016c40100000000000000000000000000000000000000040018c40100000000000000000000000000000000000000040018c4010000000000000000000000000000000000000004001ac4010000000000000000000000000000000000000004001ac40100000000000000000000000000000000000000040024c40100000000000000000000000000000000000000040026c4010000000000000000000000000000000000000004002ec4010000000000000000000000000000000000000004002ec40100000000000000000000000000000000000000040034c40100000000000000000000000000000000000000040034c40100000000000000000000000000000000000000040036c40100000000000000000000000000000000000000040036c4010000000000000000000000000092430000000004003cc4010000000000000000000000000000000000000004004ac4010000000000000000000000000000000000000004004ac4010000000000000000000000000000000000000004004cc4010000000000000000000000000000000000000004004cc40100000000000000000000000000a04300000000040052c40100000000000000000000000000000000000000040062c40100000000000000000000000000000000000000040062c40100000000000000000000000000000000000000040066c40100000000000000000000000000000000000000040066c4010000000000000000000000000000000000000004006ec40100000000000000000000000000000000000000040072c40100000000000000000000000000000000000000040072c40100000000000000000000000000ae4300000200040072c40100000000007000000000000000000000000000040072c40100000000000000000000000000000000000000040072c40100000000000000000000000000000000000000040072c40100000000000000000000000000000000000000040074c40100000000000000000000000000000000000000040076c40100000000000000000000000000000000000000040078c40100000000000000000000000000000000000000040078c40100000000000000000000000000000000000000040080c40100000000000000000000000000000000000000040080c40100000000000000000000000000000000000000040088c40100000000000000000000000000000000000000040088c4010000000000000000000000000000000000000004008ac4010000000000000000000000000000000000000004008ac4010000000000000000000000000000000000000004008ec4010000000000000000000000000000000000000004008ec40100000000000000000000000000000000000000040096c40100000000000000000000000000000000000000040098c40100000000000000000000000000000000000000040098c401000000000000000000000000000000000000000400a0c401000000000000000000000000000000000000000400a0c401000000000000000000000000000000000000000400a4c401000000000000000000000000000000000000000400a4c401000000000000000000000000000000000000000400aec401000000000000000000000000000000000000000400aec401000000000000000000000000000000000000000400b8c401000000000000000000000000000e44000000000400b8c401000000000000000000000000000000000000000400b8c401000000000000000000000000000000000000000400cec401000000000000000000000000000000000000000400cec401000000000000000000000000000000000000000400d0c401000000000000000000000000000000000000000400d4c401000000000000000000000000000000000000000400d4c401000000000000000000000000000000000000000400e2c401000000000000000000000000000000000000000400e2c401000000000000000000000000000000000000000400e2c401000000000000000000000000000000000000000400e2c401000000000000000000000000000000000000000400e4c401000000000000000000000000000000000000000400eec401000000000000000000000000001c4400000200040034c50100000000007e00000000000000000000000000040034c50100000000000000000000000000000000000000040034c50100000000000000000000000000000000000000040036c5010000000000000000000000000000000000000004003cc501000000000000000000000000000000000000000400b2c501000000000000000000000000000000000000000400b2c501000000000000000000000000000000000000000400b4c501000000000000000000000000000000000000000400bcc50100000000000000000000000000000000000000040014c60100000000000000000000000000764400000200040014c60100000000003600000000000000000000000000040014c6010000000000000000000000000000000000000004004ac60100000000000000000000000000be440000020004004ac6010000000000300000000000000000000000000004004ac6010000000000000000000000000000000000000004007ac6010000000000000000000000000000000000000004007ac6010000000000000000000000000000000000000004007cc60100000000000000000000000000000000000000040080c601000000000000000000000000000000000000000400c8c601000000000000000000000000000645000002000400c8c601000000000086000000000000000000000000000400c8c601000000000000000000000000000000000000000400cac601000000000000000000000000000000000000000400d6c601000000000000000000000000006545000000000400e4c601000000000000000000000000007345000001000100e60501000000000001000000000000009f45000000000400fec60100000000000000000000000000ad450000000004002ec70100000000000000000000000000bb450000010001002d06010000000000010000000000000000000000000004004ec70100000000000000000000000000e7450000020004004ec7010000000000680000000000000000000000000004004ec70100000000000000000000000000000000000000040050c7010000000000000000000000000000000000000004005ac701000000000000000000000000002846000002000400b6c70100000000007e000000000000000000000000000400b6c701000000000000000000000000000000000000000400b6c701000000000000000000000000000000000000000400b8c701000000000000000000000000000000000000000400bec70100000000000000000000000000824600000200040034c80100000000005200000000000000000000000000040034c80100000000000000000000000000000000000000040034c80100000000000000000000000000000000000000040036c8010000000000000000000000000000000000000004003cc80100000000000000000000000000000000000000040086c80100000000000000000000000000000000000000040086c80100000000000000000000000000000000000000040088c8010000000000000000000000000000000000000004008cc801000000000000000000000000000000000000000400dcc80100000000000000000000000000b546000002000400dcc801000000000082010000000000000000000000000400dcc801000000000000000000000000000000000000000400dec801000000000000000000000000000000000000000400ecc80100000000000000000000000000e646000000000400bec90100000000000000000000000000f44600000100010000080100000000001c00000000000000fe46000000000400c8c901000000000000000000000000000c47000000000400d2c901000000000000000000000000001a47000000000400e6c901000000000000000000000000002847000000000400eec901000000000000000000000000003647000001000100880701000000000020000000000000006047000000000400fcc901000000000000000000000000006e4700000100010066080100000000002f0000000000000099470000000004000aca0100000000000000000000000000a74700000100010095080100000000003200000000000000d24700000000040024ca0100000000000000000000000000e0470000000004002cca0100000000000000000000000000ee47000001000100e0070100000000002000000000000000184800000000040046ca010000000000000000000000000026480000010001001c080100000000001c00000000000000514800000000040050ca01000000000000000000000000005f4800000100010038080100000000002e0000000000000000000000000004005eca01000000000000000000000000008a480000020004005eca010000000000280000000000000000000000000004005eca0100000000000000000000000000e54800000000040064ca0100000000000000000000000000f348000001000100d00d01000000000050000000000000005d490000000004006eca01000000000000000000000000006b49000001000100200e0100000000005000000000000000000000000000040086ca0100000000000000000000000000000000000000040086ca0100000000000000000000000000000000000000040088ca0100000000000000000000000000d949000000000400a8ca0100000000000000000000000000e749000000000400b4ca0100000000000000000000000000f549000001000100a80701000000000018000000000000001f4a000000000400bcca01000000000000000000000000002d4a000001000100c0070100000000002000000000000000574a000000000400d2ca0100000000000000000000000000654a000001000100c70801000000000026000000000000000000000000000400e8ca0100000000000000000000000000904a000002000400e8ca01000000000068000000000000000000000000000400e8ca01000000000000000000000000000000000000000400eaca01000000000000000000000000000000000000000400eeca0100000000000000000000000000cf4a0000000004001acb0100000000000000000000000000dd4a00000000040022cb0100000000000000000000000000eb4a0000000004003ccb0100000000000000000000000000f94a000001000100ed080100000000000d00000000000000000000000000040050cb0100000000000000000000000000000000000000040050cb0100000000000000000000000000000000000000040052cb0100000000000000000000000000000000000000040054cb0100000000000000000000000000244b0000000004006ccb0100000000000000000000000000324b000001000100fa080100000000000e00000000000000000000000000040080cb0100000000000000000000000000000000000000040080cb0100000000000000000000000000000000000000040082cb0100000000000000000000000000000000000000040094cb01000000000000000000000000005d4b00000000040010cc01000000000000000000000000006b4b0000000004009ecc0100000000000000000000000000794b000000000400a8cc0100000000000000000000000000874b000000000400b2cc0100000000000000000000000000954b000000000400bccc0100000000000000000000000000a34b000000000400c6cc0100000000000000000000000000b14b000000000400d0cc01000000000000000000000000000000000000000400e6cc01000000000000000000000000000000000000000400e6cc01000000000000000000000000000000000000000400e8cc01000000000000000000000000000000000000000400eccc0100000000000000000000000000bf4b00000000040034cd010000000000000000000000000000000000000004004acd010000000000000000000000000000000000000004004acd010000000000000000000000000000000000000004004ccd0100000000000000000000000000000000000000040052cd0100000000000000000000000000cd4b0000000004008ccd0100000000000000000000000000db4b00000000040094cd0100000000000000000000000000e94b000000000400aecd0100000000000000000000000000f74b00000100010008090100000000000e000000000000000000000000000400c2cd01000000000000000000000000000000000000000400c2cd01000000000000000000000000000000000000000400c4cd01000000000000000000000000000000000000000400cacd0100000000000000000000000000224c0000000004000ace0100000000000000000000000000304c00000000040012ce01000000000000000000000000003e4c0000000004002cce01000000000000000000000000004c4c00000100010024090100000000000d00000000000000000000000000040040ce0100000000000000000000000000000000000000040040ce0100000000000000000000000000000000000000040042ce010000000000000000000000000000000000000004004ace0100000000000000000000000000774c000000000400acce0100000000000000000000000000854c000000000400b4ce0100000000000000000000000000934c000000000400cece0100000000000000000000000000a14c000001000100310901000000000012000000000000000000000000000400e2ce0100000000000000000000000000cc4c000002000400e2ce0100000000007a000000000000000000000000000400e2ce01000000000000000000000000000000000000000400e4ce01000000000000000000000000000000000000000400eace0100000000000000000000000000304d0000000004003acf010000000000000000000000000000000000000004005ccf010000000000000000000000000000000000000004005ccf010000000000000000000000000000000000000004005ecf010000000000000000000000000000000000000004006acf01000000000000000000000000003e4d000000000400c4cf01000000000000000000000000004c4d00000100010048090100000000002000000000000000000000000000040016d00100000000000000000000000000774d00000200040016d00100000000001000000000000000000000000000040016d00100000000000000000000000000000000000000040026d00100000000000000000000000000c84d00000200040026d00100000000008c00000000000000000000000000040026d00100000000000000000000000000000000000000040028d00100000000000000000000000000000000000000040030d001000000000000000000000000000000000000000400b2d001000000000000000000000000000b4e000002000400b2d00100000000004a000000000000000000000000000400b2d001000000000000000000000000000000000000000400fcd001000000000000000000000000006f4e000002000400fcd001000000000072000000000000000000000000000400fcd001000000000000000000000000000000000000000400fed00100000000000000000000000000000000000000040006d10100000000000000000000000000f04e00000000040050d10100000000000000000000000000fe4e000001000100100a0100000000001c0000000000000000000000000004006ed1010000000000000000000000000000000000000004006ed10100000000000000000000000000084f0000000004000ed20100000000000000000000000000164f00000000040024d2010000000000000000000000000000000000000004002ed20100000000000000000000000000244f0000020004002ed2010000000000280000000000000000000000000004002ed20100000000000000000000000000000000000000040030d20100000000000000000000000000000000000000040032d20100000000000000000000000000000000000000040056d20100000000000000000000000000694f00000200040056d20100000000002800000000000000000000000000040056d20100000000000000000000000000000000000000040058d2010000000000000000000000000000000000000004005ad2010000000000000000000000000000000000000004007ed20100000000000000000000000000ae4f0000020004007ed2010000000000140100000000000000000000000004007ed20100000000000000000000000000000000000000040080d20100000000000000000000000000000000000000040098d20100000000000000000000000000000000000000040092d30100000000000000000000000000c95000000200040092d30100000000006c00000000000000000000000000040092d301000000000000000000000000000000000000000400fed301000000000000000000000000006e51000002000400fed30100000000007e030000000000000000000000000400fed30100000000000000000000000000000000000000040000d4010000000000000000000000000000000000000004001ad40100000000000000000000000000bc5200000200040082da010000000000e8020000000000002c530000020004007cd7010000000000060300000000000093530000020004006add010000000000d002000000000000f9530000020004003ae0010000000000ae0200000000000000000000000004007cd7010000000000000000000000000000000000000004007cd7010000000000000000000000000000000000000004007ed70100000000000000000000000000000000000000040098d7010000000000000000000000000057540000000004003eda010000000000000000000000000065540000010001009e0b0100000000001b0000000000000090540000000004004ada01000000000000000000000000009e5400000000040058da0100000000000000000000000000ac5400000000040062da0100000000000000000000000000ba540000000004006cda0100000000000000000000000000000000000000040082da0100000000000000000000000000000000000000040082da0100000000000000000000000000000000000000040084da010000000000000000000000000000000000000004009eda0100000000000000000000000000c85400000000040046dd0100000000000000000000000000d65400000000040054dd010000000000000000000000000000000000000004006add010000000000000000000000000000000000000004006add010000000000000000000000000000000000000004006cdd0100000000000000000000000000000000000000040086dd0100000000000000000000000000e454000000000400f2df0100000000000000000000000000f254000000000400fedf010000000000000000000000000000550000000004000ce001000000000000000000000000000e550000000004001ae001000000000000000000000000001c5500000000040024e0010000000000000000000000000000000000000004003ae0010000000000000000000000000000000000000004003ae0010000000000000000000000000000000000000004003ce00100000000000000000000000000000000000000040056e001000000000000000000000000002a55000000000400d2e201000000000000000000000000000000000000000400e8e201000000000000000000000000003855000002000400e8e201000000000028000000000000000000000000000400e8e201000000000000000000000000000000000000000400eae201000000000000000000000000000000000000000400ece20100000000000000000000000000000000000000040010e301000000000000000000000000007d5500000200040010e30100000000002800000000000000000000000000040010e30100000000000000000000000000000000000000040012e30100000000000000000000000000000000000000040014e30100000000000000000000000000000000000000040038e30100000000000000000000000000c25500000200040038e30100000000002801000000000000000000000000040038e3010000000000000000000000000000000000000004003ae30100000000000000000000000000000000000000040050e30100000000000000000000000000000000000000040060e40100000000000000000000000000dd5600000200040060e40100000000006800000000000000000000000000040060e40100000000000000000000000000000000000000040062e40100000000000000000000000000000000000000040070e401000000000000000000000000000000000000000400c8e401000000000000000000000000008257000002000400c8e401000000000004030000000000000000000000000400c8e401000000000000000000000000000000000000000400cce40100000000000000000000000000000000000000040000e50100000000000000000000000000d058000002000400cce701000000000066000000000000009859000002000400f8ea0100000000004602000000000000085a00000200040032e8010000000000c6020000000000006f5a0000020004003eed0100000000008e02000000000000d55a000002000400ccef01000000000002020000000000000000000000000400cce701000000000000000000000000000000000000000400cce70100000000000000000000000000000000000000040032e80100000000000000000000000000000000000000040032e80100000000000000000000000000000000000000040036e8010000000000000000000000000000000000000004006ae80100000000000000000000000000335b000000000400b4ea0100000000000000000000000000415b000000000400c0ea01000000000000000000000000004f5b000000000400ceea01000000000000000000000000005d5b000000000400d8ea01000000000000000000000000006b5b000000000400e2ea01000000000000000000000000000000000000000400f8ea01000000000000000000000000000000000000000400f8ea01000000000000000000000000000000000000000400faea0100000000000000000000000000000000000000040014eb0100000000000000000000000000795b0000000004001aed0100000000000000000000000000875b00000000040028ed010000000000000000000000000000000000000004003eed010000000000000000000000000000000000000004003eed0100000000000000000000000000000000000000040042ed0100000000000000000000000000000000000000040076ed0100000000000000000000000000955b00000000040084ef0100000000000000000000000000a35b00000000040090ef0100000000000000000000000000b15b0000000004009eef0100000000000000000000000000bf5b000000000400acef0100000000000000000000000000cd5b000000000400b6ef01000000000000000000000000000000000000000400ccef01000000000000000000000000000000000000000400ccef01000000000000000000000000000000000000000400ceef01000000000000000000000000000000000000000400e8ef0100000000000000000000000000db5b000000000400b8f101000000000000000000000000000000000000000400cef10100000000000000000000000000e95b000002000400cef101000000000036290000000000000000000000000400cef101000000000000000000000000000000000000000400d2f101000000000000000000000000000000000000000400fcf10100000000000000000000000000195c000002000400a82002000000000006040000000000005c5c000002000400962e0200000000005001000000000000945c000002000400e62f0200000000000c03000000000000d45c000002000400ae24020000000000e8090000000000000000000000000400041b0200000000000000000000000000055d000000000500b0c90200000000000000000000000000105d000002000400041b0200000000008e000000000000000000000000000400041b02000000000000000000000000000000000000000400061b020000000000000000000000000000000000000004000c1b02000000000000000000000000005d5d000000000400261b02000000000000000000000000000000000000000400921b02000000000000000000000000006b5d000002000400921b020000000000cc010000000000000000000000000400921b02000000000000000000000000000000000000000400961b02000000000000000000000000000000000000000400ae1b0200000000000000000000000000a35d000000000400c81b0200000000000000000000000000b15d000002000400ba360200000000006a00000000000000df5d0000020004005e1d020000000000f600000000000000225e000000000400b81c0200000000000000000000000000305e000000000400dc1c02000000000000000000000000003e5e000002000400541e020000000000540200000000000000000000000004005e1d020000000000000000000000000000000000000004005e1d02000000000000000000000000000000000000000400621d02000000000000000000000000000000000000000400761d02000000000000000000000000000000000000000400541e02000000000000000000000000000000000000000400541e02000000000000000000000000000000000000000400581e02000000000000000000000000000000000000000400701e02000000000000000000000000000000000000000400a82002000000000000000000000000000000000000000400a82002000000000000000000000000000000000000000400aa2002000000000000000000000000000000000000000400c0200200000000000000000000000000815e000000000400982402000000000000000000000000008f5e000001000100300a0100000000002e000000000000000000000000000400ae2402000000000000000000000000000000000000000400ae2402000000000000000000000000000000000000000400b02402000000000000000000000000000000000000000400c82402000000000000000000000000000000000000000400962e0200000000000000000000000000ba5e000000000500b8c90200000000000000000000000000c55e000000000500c0c90200000000000000000000000000d05e000000000500c8c90200000000000000000000000000db5e000000000500d0c902000000000000000000000000000000000000000400962e02000000000000000000000000000000000000000400982e02000000000000000000000000000000000000000400aa2e0200000000000000000000000000e65e000000000400d62e0200000000000000000000000000f45e000000000400de2e0200000000000000000000000000025f000000000400f82e0200000000000000000000000000105f000000000400002f02000000000000000000000000001e5f000000000400d22f02000000000000000000000000000000000000000400e62f02000000000000000000000000000000000000000400e62f02000000000000000000000000000000000000000400e82f02000000000000000000000000000000000000000400023002000000000000000000000000002c5f000002000400f232020000000000c8030000000000000000000000000400f23202000000000000000000000000000000000000000400f23202000000000000000000000000000000000000000400f43202000000000000000000000000000000000000000400043302000000000000000000000000000000000000000400ba3602000000000000000000000000000000000000000400ba3602000000000000000000000000000000000000000400bc3602000000000000000000000000000000000000000400c4360200000000000000000000000000705f000000000400ec3602000000000000000000000000000000000000000400243702000000000000000000000000007e5f000000000500d8c90200000000000000000000000000895f00000200040024370200000000008e0000000000000000000000000004002437020000000000000000000000000000000000000004002637020000000000000000000000000000000000000004002c370200000000000000000000000000d65f000000000400463702000000000000000000000000000000000000000400b2370200000000000000000000000000e45f000002000400b23702000000000072000000000000000000000000000400b23702000000000000000000000000000000000000000400b43702000000000000000000000000000000000000000400bc3702000000000000000000000000006560000000000400103802000000000000000000000000000000000000000400243802000000000000000000000000000000000000000400243802000000000000000000000000007360000000000400263802000000000000000000000000008160000000000100880101000000000000000000000000008c6000000000040036380200000000000000000000000000966000000000040038380200000000000000000000000000a0600000000004003a380200000000000000000000000000aa600000000004003e380200000000000000000000000000b4600000000004004238020000000000000000000000000000000000000004004c38020000000000000000000000000000000000000004004c38020000000000000000000000000000000000000004006838020000000000000000000000000000000000000004006838020000000000000000000000000000000000000004006c380200000000000000000000000000000000000000040084380200000000000000000000000000be60000000000400ba380200000000000000000000000000000000000000040042390200000000000000000000000000000000000000040042390200000000000000000000000000000000000000040044390200000000000000000000000000000000000000040050390200000000000000000000000000cc600000020004006c3b02000000000032000000000000003e610000000004004c3b02000000000000000000000000004c61000000000400543b02000000000000000000000000005a61000001000100900a010000000000200000000000000000000000000004006c3b020000000000000000000000000000000000000004006c3b020000000000000000000000000000000000000004006e3b02000000000000000000000000000000000000000400723b020000000000000000000000000000000000000004009e3b020000000000000000000000000000000000000004009e3b02000000000000000000000000000000000000000400a03b02000000000000000000000000000000000000000400b63b02000000000000000000000000008561000000000400743e02000000000000000000000000009361000000000400883e0200000000000000000000000000a161000001000100500d0100000000002b00000000000000cd61000000000400963e0200000000000000000000000000db610000000004009e3e02000000000000000000000000000000000000000400b63e02000000000000000000000000000000000000000400b63e02000000000000000000000000000000000000000400b83e02000000000000000000000000000000000000000400d23e0200000000000000000000000000e96100000000040000420200000000000000000000000000f7610000000004001442020000000000000000000000000005620000000004001c4202000000000000000000000000001362000001000100b00a01000000000020000000000000003e62000000000400344202000000000000000000000000004c620000010001007b0d010000000000290000000000000000000000000004004242020000000000000000000000000000000000000004004242020000000000000000000000000000000000000004004442020000000000000000000000000000000000000004005e4202000000000000000000000000007862000000000400904502000000000000000000000000008662000000000400a44502000000000000000000000000009462000000000400ac450200000000000000000000000000a262000000000400c4450200000000000000000000000000b062000001000100a40d0100000000002c000000000000000000000000000400d24502000000000000000000000000000000000000000400d24502000000000000000000000000000000000000000400d44502000000000000000000000000000000000000000400ee450200000000000000000000000000dc620000000004009e490200000000000000000000000000ea62000000000400b2490200000000000000000000000000f862000000000400ba4902000000000000000000000000000663000000000400ca4902000000000000000000000000001463000000000400d24902000000000000000000000000002263000000000400e24902000000000000000000000000003063000000000400ea4902000000000000000000000000003e63000000000400f44902000000000000000000000000004c63000000000400fc4902000000000000000000000000000000000000000400204a02000000000000000000000000000000000000000400204a02000000000000000000000000000000000000000400224a020000000000000000000000000000000000000004002e4a02000000000000000000000000005a63000000000400804b02000000000000000000000000000000000000000400a64b02000000000000000000000000006863000002000400a64b02000000000056020000000000000000000000000400a64b02000000000000000000000000000000000000000400a84b02000000000000000000000000000000000000000400c24b0200000000000000000000000000a863000000000400c84d0200000000000000000000000000b663000000000400dc4d0200000000000000000000000000c463000000000400e44d02000000000000000000000000000000000000000400fc4d02000000000000000000000000000000000000000400fc4d02000000000000000000000000000000000000000400fe4d02000000000000000000000000000000000000000400064e0200000000000000000000000000d263000000000400744e0200000000000000000000000000e0630000000004007c4e02000000000000000000000000000000000000000400964e02000000000000000000000000000000000000000400964e02000000000000000000000000000000000000000400984e020000000000000000000000000000000000000004009e4e0200000000000000000000000000ee63000000000400964f0200000000000000000000000000fc630000000004009e4f02000000000000000000000000000a64000000000400a84f02000000000000000000000000001864000000000400b04f02000000000000000000000000002664000000000400c04f02000000000000000000000000003464000000000400c84f02000000000000000000000000004264000000000400d84f02000000000000000000000000005064000000000400e04f02000000000000000000000000005e64000000000400fa4f02000000000000000000000000006c6400000100010016090100000000000e0000000000000000000000000004000e50020000000000000000000000000000000000000004000e50020000000000000000000000000000000000000004001050020000000000000000000000000000000000000004002a500200000000000000000000000000976400000000040020520200000000000000000000000000a56400000000040034520200000000000000000000000000b3640000000004003c520200000000000000000000000000c1640000000004005452020000000000000000000000000000000000000004006252020000000000000000000000000000000000000004006252020000000000000000000000000000000000000004006652020000000000000000000000000000000000000004009a520200000000000000000000000000cf64000000000400c8580200000000000000000000000000dd640000000004008a590200000000000000000000000000eb6400000100010080020100000000001c00000000000000f164000000000400b4590200000000000000000000000000ff64000000000400bc5902000000000000000000000000000d65000001000100d00a01000000000020000000000000000000000000000400d45902000000000000000000000000000000000000000400d45902000000000000000000000000000000000000000400d85902000000000000000000000000000000000000000400e45902000000000000000000000000000000000000000400485a02000000000000000000000000000000000000000400485a020000000000000000000000000000000000000004004c5a02000000000000000000000000000000000000000400805a02000000000000000000000000000000000000000400805a02000000000000000000000000000000000000000400825a02000000000000000000000000003865000000000400dc5b02000000000000000000000000004665000000000400967502000000000000000000000000005465000000000400b87502000000000000000000000000006265000000000400228802000000000000000000000000007065000000000100b00101000000000000000000000000007b650000000004000093020000000000000000000000000087650000000004005688020000000000000000000000000093650000000004002a8a02000000000000000000000000009f650000000004008e8c0200000000000000000000000000ab650000000004004a8e0200000000000000000000000000b7650000000004009a8e0200000000000000000000000000c36500000000040018930200000000000000000000000000d1650000000004002a930200000000000000000000000000df6500000000040038930200000000000000000000000000ed6500000000040046930200000000000000000000000000fb650000000004005093020000000000000000000000000009660000000004005a93020000000000000000000000000017660000000004006493020000000000000000000000000025660000000004007e93020000000000000000000000000033660000000004009493020000000000000000000000000041660000000004009e9302000000000000000000000000004f66000000000400ac9302000000000000000000000000005d66000000000400c09302000000000000000000000000006b66000000000400ca9302000000000000000000000000007966000000000400d49302000000000000000000000000008766000000000400de9302000000000000000000000000009566000000000400e8930200000000000000000000000000a366000000000400f2930200000000000000000000000000b16600000000040006940200000000000000000000000000bf6600000000040010940200000000000000000000000000cd660000000004001a940200000000000000000000000000db6600000000040024940200000000000000000000000000e9660000000004002e940200000000000000000000000000f7660000000004003894020000000000000000000000000005670000000004005a94020000000000000000000000000013670000000004006494020000000000000000000000000021670000000004006e9402000000000000000000000000002f670000000004007e9402000000000000000000000000003d67000000000400889402000000000000000000000000000000000000000400929402000000000000000000000000004b67000001000800a0ca02000000000000100800000000007a67000001000800a0da0a00000000000010000000000000af67000001000100dc030100000000002300000000000000da6700000100010010040100000000003300000000000000056800000100010068090100000000000a00000000000000306800000100010072090100000000000a000000000000005b680000010001007c090100000000000b00000000000000866800000100010087090100000000000600000000000000b1680000010001008d090100000000000600000000000000dc680000010001009309010000000000090000000000000007690000010001009c0901000000000006000000000000000000000000000a00000000000000000000000000000000000000000000000d00752b00000000000000000000000000000000000000000d00604600000000000000000000000000003269000000001100000000000000000000000000000000000000000000000d002b1300000000000000000000000000000000000000000c00701100000000000000000000000000000000000000000d00742f00000000000000000000000000000000000000000d00000000000000000000000000000000000000000000000d007c4f00000000000000000000000000000000000000000d00643800000000000000000000000000000000000000000d00953f00000000000000000000000000000000000000000d00190f00000000000000000000000000000000000000000a00740000000000000000000000000000000000000000000d005a1700000000000000000000000000004669000000001100880000000000000000000000000000000000000000000c00a01100000000000000000000000000000000000000000d003b1a00000000000000000000000000000000000000000d00840500000000000000000000000000000000000000000d002f0d00000000000000000000000000000000000000000d00901700000000000000000000000000000000000000000d00dc3500000000000000000000000000000000000000000d00dd0c00000000000000000000000000000000000000000d00ab3f00000000000000000000000000000000000000000d00973300000000000000000000000000000000000000000d00e63800000000000000000000000000000000000000000d00182500000000000000000000000000000000000000000d009a2a00000000000000000000000000000000000000000d006c2300000000000000000000000000000000000000000d00eb2c00000000000000000000000000000000000000000d00d14900000000000000000000000000000000000000000d00ba3b00000000000000000000000000000000000000000d006f3a00000000000000000000000000000000000000000d00770c00000000000000000000000000000000000000000d00f90300000000000000000000000000000000000000000d005f0d00000000000000000000000000000000000000000d00ae4200000000000000000000000000000000000000000d00b03300000000000000000000000000000000000000000d008d1800000000000000000000000000000000000000000d00ff0b00000000000000000000000000000000000000000d00d53700000000000000000000000000000000000000000d00a60000000000000000000000000000000000000000000d00794a00000000000000000000000000000000000000000d00fd1300000000000000000000000000000000000000000d00574400000000000000000000000000000000000000000d00244900000000000000000000000000000000000000000d00900500000000000000000000000000000000000000000d00b80800000000000000000000000000000000000000000d00cc0000000000000000000000000000000000000000000d000b2a00000000000000000000000000000000000000000d00933300000000000000000000000000000000000000000d005b1300000000000000000000000000000000000000000d00903400000000000000000000000000000000000000000d00fd4b00000000000000000000000000000000000000000d00542900000000000000000000000000000000000000000d007b4100000000000000000000000000000000000000000d00361400000000000000000000000000000000000000000d00c84900000000000000000000000000000000000000000d008f3e00000000000000000000000000000000000000000d00544c00000000000000000000000000000000000000000d004f3100000000000000000000000000000000000000000d00fc1600000000000000000000000000000000000000000d00763800000000000000000000000000000000000000000c00000000000000000000000000000000000000000000000c00400000000000000000000000000000000000000000000c00700000000000000000000000000000000000000000000c00a00000000000000000000000000000000000000000000d00550c00000000000000000000000000000000000000000d00472d00000000000000000000000000000000000000000d00c03e00000000000000000000000000000000000000000d00441b00000000000000000000000000000000000000000d00f20400000000000000000000000000000000000000000d00c11600000000000000000000000000000000000000000d00b41000000000000000000000000000000000000000000d00aa3000000000000000000000000000000000000000000d004e2b00000000000000000000000000000000000000000d002a2b00000000000000000000000000000000000000000d00011500000000000000000000000000000000000000000d00581d00000000000000000000000000000000000000000d008b4700000000000000000000000000000000000000000d00c54a00000000000000000000000000000000000000000d001d3c00000000000000000000000000000000000000000d00761500000000000000000000000000000000000000000d00ef3000000000000000000000000000000000000000000c00200900000000000000000000000000000000000000000c00500900000000000000000000000000000000000000000c00800900000000000000000000000000000000000000000c00b00900000000000000000000000000000000000000000c00e00900000000000000000000000000000000000000000d00c60700000000000000000000000000000000000000000d00733500000000000000000000000000000000000000000d000f0f00000000000000000000000000000000000000000d00f52800000000000000000000000000000000000000000c00100e00000000000000000000000000000000000000000c00400e00000000000000000000000000000000000000000c00700e00000000000000000000000000000000000000000c00a00e00000000000000000000000000000000000000000c00d00e00000000000000000000000000000000000000000d004b4800000000000000000000000000000000000000000d00af4800000000000000000000000000000000000000000c00000f00000000000000000000000000000000000000000c00300f00000000000000000000000000000000000000000c00600f00000000000000000000000000000000000000000c00900f00000000000000000000000000000000000000000c00c00f00000000000000000000000000000000000000000d00210800000000000000000000000000000000000000000d001f0300000000000000000000000000000000000000000c00801000000000000000000000000000000000000000000c00b01000000000000000000000000000000000000000000c00e01000000000000000000000000000000000000000000c00101100000000000000000000000000000000000000000c00401100000000000000000000000000000000000000000d00d74d00000000000000000000000000000000000000000d00e90a00000000000000000000000000000000000000000d001e0b00000000000000000000000000000000000000000d007f0300000000000000000000000000000000000000000d00533100000000000000000000000000000000000000000d00c94c00000000000000000000000000000000000000000d00434400000000000000000000000000000000000000000d006b0d00000000000000000000000000000000000000000d00880500000000000000000000000000000000000000000d00890200000000000000000000000000000000000000000d00cc3400000000000000000000000000000000000000000c00d00000000000000000000000000000000000000000000c00100100000000000000000000000000000000000000000c00400100000000000000000000000000000000000000000c00700100000000000000000000000000000000000000000c00a00100000000000000000000000000000000000000000c00d00100000000000000000000000000000000000000000c00000200000000000000000000000000000000000000000c00300200000000000000000000000000000000000000000c00800200000000000000000000000000000000000000000d00784b00000000000000000000000000000000000000000d00e53000000000000000000000000000000000000000000c00b00200000000000000000000000000000000000000000c00e00200000000000000000000000000000000000000000c00100300000000000000000000000000000000000000000c00400300000000000000000000000000000000000000000c00700300000000000000000000000000000000000000000c00a00300000000000000000000000000000000000000000c00d00300000000000000000000000000000000000000000c00000400000000000000000000000000000000000000000c00300400000000000000000000000000000000000000000c00800400000000000000000000000000000000000000000c00b00400000000000000000000000000000000000000000c00000500000000000000000000000000000000000000000c00300500000000000000000000000000000000000000000c00800500000000000000000000000000000000000000000c00b00500000000000000000000000000000000000000000c00f00500000000000000000000000000000000000000000c00600600000000000000000000000000000000000000000c00b00600000000000000000000000000000000000000000c00f00600000000000000000000000000000000000000000c00200700000000000000000000000000000000000000000c00500700000000000000000000000000000000000000000d008b3b00000000000000000000000000000000000000000d00043000000000000000000000000000000000000000000d00981800000000000000000000000000000000000000000d003d2d00000000000000000000000000000000000000000d00123400000000000000000000000000000000000000000d001d2b00000000000000000000000000000000000000000d00c12800000000000000000000000000000000000000000d00ea1d00000000000000000000000000000000000000000d00db0700000000000000000000000000000000000000000d00fe2400000000000000000000000000000000000000000d00c51b00000000000000000000000000000000000000000d00591800000000000000000000000000000000000000000d00e73100000000000000000000000000000000000000000d00ed3100000000000000000000000000000000000000000d00874d00000000000000000000000000000000000000000d007f1b00000000000000000000000000000000000000000d00ac0900000000000000000000000000000000000000000d00434d00000000000000000000000000000000000000000d00171000000000000000000000000000000000000000000d00d10900000000000000000000000000000000000000000d00943c00000000000000000000000000000000000000000c00800700000000000000000000000000000000000000000c00b00700000000000000000000000000000000000000000c00e00700000000000000000000000000000000000000000c00100800000000000000000000000000000000000000000c00400800000000000000000000000000000000000000000c00700800000000000000000000000000000000000000000c00a00800000000000000000000000000000000000000000c00e00800000000000000000000000000000000000000000d00f10100000000000000000000000000000000000000000d00244000000000000000000000000000000000000000000d000c3c00000000000000000000000000000000000000000d003b3b00000000000000000000000000000000000000000d007e3800000000000000000000000000000000000000000c00100a00000000000000000000000000000000000000000c00400a00000000000000000000000000000000000000000c00700a00000000000000000000000000000000000000000c00a00a00000000000000000000000000000000000000000c00d00a00000000000000000000000000000000000000000c00000b00000000000000000000000000000000000000000d00b14000000000000000000000000000000000000000000d00454800000000000000000000000000000000000000000d00920400000000000000000000000000000000000000000d003d1b00000000000000000000000000000000000000000d00a32400000000000000000000000000000000000000000d00432b00000000000000000000000000000000000000000d00474d00000000000000000000000000000000000000000d00664a00000000000000000000000000000000000000000d006f0a00000000000000000000000000000000000000000c00b00b00000000000000000000000000000000000000000c00e00b00000000000000000000000000000000000000000c00100c00000000000000000000000000000000000000000c00400c00000000000000000000000000000000000000000c00700c00000000000000000000000000000000000000000c00b00c00000000000000000000000000000000000000000d00641e00000000000000000000000000000000000000000d006d4b00000000000000000000000000000000000000000d00291e00000000000000000000000000000000000000000d000f3000000000000000000000000000000000000000000d00a30900000000000000000000000000000000000000000d000b3800000000000000000000000000000000000000000d00321b00000000000000000000000000000000000000000d00143000000000000000000000000000000000000000000d00ec0400000000000000000000000000000000000000000d00cf0e00000000000000000000000000000000000000000d00114d00000000000000000000000000000000000000000d00503000000000000000000000000000000000000000000d00dc3a00000000000000000000000000000000000000000d004b0500000000000000000000000000000000000000000c00f00c00000000000000000000000000000000000000000c00200d00000000000000000000000000000000000000000c00500d00000000000000000000000000000000000000000c00800d00000000000000000000000000000000000000000c00b00d00000000000000000000000000000000000000000c00e00d00000000000000000000000000000000000000000d00553400000000000000000000000000000000000000000d00932400000000000000000000000000000000000000000d00d43200000000000000000000000000000000000000000c00300b00000000000000000000000000000000000000000d00ae1900000000000000000000000000000000000000000d00da3200000000000000000000000000000000000000000d00144800000000000000000000000000000000000000000d00514f00000000000000000000000000000000000000000d00a74b00000000000000000000000000000000000000000d00774500000000000000000000000000000000000000000d00a24500000000000000000000000000000000000000000c00700b00000000000000000000000000000000000000000d00e53a00000000000000000000000000000000000000000d002a0a00000000000000000000000000000000000000000d00da1000000000000000000000000000000000000000000d00d30c00000000000000000000000000000000000000000d004b3300000000000000000000000000000000000000000d00251100000000000000000000000000000000000000000d00db3c00000000000000000000000000000000000000000d00ce4d00000000000000000000000000000000000000000d004d4c00000000000000000000000000000000000000000d00340a00000000000000000000000000000000000000000d00b54f00000000000000000000000000000000000000000d00242f00000000000000000000000000000000000000000d00d00700000000000000000000000000000000000000000d002a2f00000000000000000000000000000000000000000d00b01000000000000000000000000000000000000000000d00df3c00000000000000000000000000000000000000000d00ab0a00000000000000000000000000000000000000000d008e1100000000000000000000000000000000000000000d009d3400000000000000000000000000000000000000000d00a11e00000000000000000000000000000000000000000d00202500000000000000000000000000000000000000000d00663600000000000000000000000000000000000000000d000e4900000000000000000000000000000000000000000d00153e00000000000000000000000000000000000000000d00c10100000000000000000000000000000000000000000d00712c00000000000000000000000000000000000000000d00764400000000000000000000000000000000000000000d006b4e00000000000000000000000000000000000000000d005a4100000000000000000000000000000000000000000d00a01c00000000000000000000000000000000000000000d00064000000000000000000000000000000000000000000d00383900000000000000000000000000000000000000000d00120000000000000000000000000000000000000000000d00a41b00000000000000000000000000000000000000000d00812f00000000000000000000000000000000000000000d00094d00000000000000000000000000000000000000000d00e13400000000000000000000000000000000000000000d007c2300000000000000000000000000000000000000000d008c2300000000000000000000000000000000000000000d004b3700000000000000000000000000000000000000000d00614e00000000000000000000000000000000000000000d00ef3900000000000000000000000000000000000000000d00740b00000000000000000000000000000000000000000d00ff3d00000000000000000000000000000000000000000d004d0c00000000000000000000000000000000000000000d001a1d00000000000000000000000000000000000000000d002c4500000000000000000000000000000000000000000d008a1200000000000000000000000000000000000000000d00d11b00000000000000000000000000000000000000000d00501c00000000000000000000000000000000000000000d00fc2900000000000000000000000000000000000000000d00404700000000000000000000000000000000000000000d009a4a00000000000000000000000000000000000000000d002c2700000000000000000000000000000000000000000d00fb4000000000000000000000000000000000000000000d00180600000000000000000000000000000000000000000d00124100000000000000000000000000000000000000000d00924400000000000000000000000000000000000000000d00620900000000000000000000000000000000000000000d003a2a00000000000000000000000000000000000000000d00862a00000000000000000000000000000000000000000d00443b00000000000000000000000000000000000000000d00ee3d00000000000000000000000000000000000000000d00b41a00000000000000000000000000000000000000000d00d11200000000000000000000000000000000000000000d00e64400000000000000000000000000000000000000000d002f3200000000000000000000000000000000000000000d00c62700000000000000000000000000000000000000000d00da0900000000000000000000000000000000000000000d005b0e00000000000000000000000000000000000000000d002b1900000000000000000000000000000000000000000d004c0400000000000000000000000000000000000000000d000a1b00000000000000000000000000000000000000000d00b60700000000000000000000000000000000000000000d00fa4500000000000000000000000000000000000000000d00c93c00000000000000000000000000000000000000000d00b40300000000000000000000000000000000000000000d00af0500000000000000000000000000000000000000000d00d93400000000000000000000000000000000000000000d00613700000000000000000000000000000000000000000d00f62a00000000000000000000000000000000000000000d00f20d00000000000000000000000000000000000000000d00ff1200000000000000000000000000000000000000000d00844100000000000000000000000000000000000000000d00fe3300000000000000000000000000000000000000000d00793a00000000000000000000000000000000000000000d00fa0100000000000000000000000000000000000000000d00ee4900000000000000000000000000000000000000000d00403200000000000000000000000000000000000000000d00cd1800000000000000000000000000000000000000000d00e91500000000000000000000000000000000000000000d009e0d00000000000000000000000000000000000000000d00801500000000000000000000000000000000000000000d00e73e00000000000000000000000000000000000000000d005e1d00000000000000000000000000000000000000000d00a64000000000000000000000000000000000000000000d00083000000000000000000000000000000000000000000d00391900000000000000000000000000000000000000000d00f53e00000000000000000000000000000000000000000d002d3f00000000000000000000000000000000000000000d002c4b00000000000000000000000000000000000000000d00db1d00000000000000000000000000000000000000000d00721000000000000000000000000000000000000000000d00f84100000000000000000000000000000000000000000d007a2f00000000000000000000000000000000000000000d00b62b00000000000000000000000000000000000000000d00984600000000000000000000000000000000000000000d005e1300000000000000000000000000000000000000000d002b2500000000000000000000000000000000000000000d00b53f00000000000000000000000000000000000000000d00fc4200000000000000000000000000000000000000000d007b3900000000000000000000000000000000000000000d00f60000000000000000000000000000000000000000000d00ec0800000000000000000000000000000000000000000d00b60f00000000000000000000000000000000000000000d00a61100000000000000000000000000000000000000000d00ac1100000000000000000000000000000000000000000d00602900000000000000000000000000000000000000000d00ea3c00000000000000000000000000000000000000000d00670d00000000000000000000000000000000000000000d00cf4300000000000000000000000000000000000000000d00b61100000000000000000000000000000000000000000d00704a00000000000000000000000000000000000000000d005d3100000000000000000000000000000000000000000d00613100000000000000000000000000000000000000000d00a61e00000000000000000000000000000000000000000d00e84d00000000000000000000000000000000000000000d00ad4600000000000000000000000000000000000000000d00c32000000000000000000000000000000000000000000d00e14d00000000000000000000000000000000000000000d002b0800000000000000000000000000000000000000000d009e1300000000000000000000000000000000000000000d000c0000000000000000000000000000000000000000000d00174900000000000000000000000000000000000000000d00a51700000000000000000000000000000000000000000d00590000000000000000000000000000000000000000000d00961c00000000000000000000000000000000000000000d00630600000000000000000000000000000000000000000d00822700000000000000000000000000000000000000000d006c1400000000000000000000000000000000000000000d00d32300000000000000000000000000000000000000000d00df0800000000000000000000000000000000000000000d004b4900000000000000000000000000000000000000000d00712200000000000000000000000000000000000000000d00844a00000000000000000000000000000000000000000d00822200000000000000000000000000000000000000000d00080000000000000000000000000000000000000000000d00280b00000000000000000000000000000000000000000d008c1b00000000000000000000000000000000000000000d00230f00000000000000000000000000000000000000000d00a14600000000000000000000000000000000000000000d00652000000000000000000000000000000000000000000d002b0900000000000000000000000000000000000000000d00a51a00000000000000000000000000000000000000000d001f4100000000000000000000000000000000000000000d00231400000000000000000000000000000000000000000d002a2c00000000000000000000000000000000000000000d00d20100000000000000000000000000000000000000000d00584c00000000000000000000000000000000000000000d00f14d00000000000000000000000000000000000000000d001f0100000000000000000000000000000000000000000d00da1b00000000000000000000000000000000000000000d00bb3200000000000000000000000000000000000000000d00172800000000000000000000000000000000000000000d00620c00000000000000000000000000000000000000000d005a4500000000000000000000000000000000000000000d00e82d00000000000000000000000000000000000000000d00c93200000000000000000000000000000000000000000d00680b00000000000000000000000000000000000000000d00ba4000000000000000000000000000000000000000000d00f43f00000000000000000000000000000000000000000d00bf2b00000000000000000000000000000000000000000d00c23900000000000000000000000000000000000000000d00d80f00000000000000000000000000000000000000000d00fe2b00000000000000000000000000000000000000000d00172300000000000000000000000000000000000000000d00592300000000000000000000000000000000000000000d003d3900000000000000000000000000000000000000000d00e33600000000000000000000000000000000000000000d00b62900000000000000000000000000000000000000000d008d4a00000000000000000000000000000000000000000d00a80d00000000000000000000000000000000000000000d000e2c00000000000000000000000000000000000000000d00e93600000000000000000000000000000000000000000d00253700000000000000000000000000000000000000000d000a0400000000000000000000000000000000000000000d00964000000000000000000000000000000000000000000d00a73300000000000000000000000000000000000000000d00240100000000000000000000000000000000000000000d00ab0500000000000000000000000000000000000000000d00174b00000000000000000000000000000000000000000d00e54e00000000000000000000000000000000000000000d001f4b00000000000000000000000000000000000000000d00652800000000000000000000000000000000000000000d006a2e00000000000000000000000000000000000000000d00263500000000000000000000000000000000000000000d00204900000000000000000000000000000000000000000d00b63d00000000000000000000000000000000000000000d00b71b00000000000000000000000000000000000000000d00a33400000000000000000000000000000000000000000d00570f00000000000000000000000000000000000000000d00822d00000000000000000000000000000000000000000d006a1500000000000000000000000000000000000000000d00bd4700000000000000000000000000000000000000000d00bb4a00000000000000000000000000000000000000000d00a20d00000000000000000000000000000000000000000d00ec0000000000000000000000000000000000000000000d00401a00000000000000000000000000000000000000000d00e03600000000000000000000000000000000000000000d008a2400000000000000000000000000000000000000000d00233c00000000000000000000000000000000000000000d00342b00000000000000000000000000000000000000000d00954700000000000000000000000000000000000000000d00f63100000000000000000000000000000000000000000d006b3a00000000000000000000000000000000000000000d001a4d00000000000000000000000000000000000000000d001f2c00000000000000000000000000000000000000000d007e0900000000000000000000000000000000000000000d00e50800000000000000000000000000000000000000000d00a03300000000000000000000000000000000000000000d00790f00000000000000000000000000000000000000000d009c0500000000000000000000000000000000000000000d00034700000000000000000000000000000000000000000d00df3d00000000000000000000000000000000000000000d00ba0300000000000000000000000000000000000000000d00824400000000000000000000000000000000000000000d00f60600000000000000000000000000000000000000000d00a70e00000000000000000000000000000000000000000d007b4200000000000000000000000000000000000000000d00bb3c00000000000000000000000000000000000000000d00bc2f00000000000000000000000000000000000000000d00ae4a00000000000000000000000000000000000000000d001e4a00000000000000000000000000000000000000000d00444f00000000000000000000000000000000000000000d00ec2a00000000000000000000000000000000000000000d002d1700000000000000000000000000000000000000000d00e93000000000000000000000000000000000000000000d00604000000000000000000000000000000000000000000d00091300000000000000000000000000000000000000000d00411000000000000000000000000000000000000000000d004b3400000000000000000000000000000000000000000d00103300000000000000000000000000000000000000000d00644500000000000000000000000000000000000000000d00051b00000000000000000000000000000000000000000d00bc2700000000000000000000000000000000000000000d00554800000000000000000000000000000000000000000d001c3500000000000000000000000000000000000000000d00c20200000000000000000000000000000000000000000d00fa1400000000000000000000000000000000000000000d00180500000000000000000000000000000000000000000d001d1300000000000000000000000000000000000000000d00664b00000000000000000000000000000000000000000d00313500000000000000000000000000000000000000000d00e11900000000000000000000000000000000000000000d00320700000000000000000000000000000000000000000d00823a00000000000000000000000000000000000000000d00740700000000000000000000000000000000000000000d003a3f00000000000000000000000000000000000000000d00063300000000000000000000000000000000000000000d000b4200000000000000000000000000000000000000000d000d0a00000000000000000000000000000000000000000d00112800000000000000000000000000000000000000000d00211900000000000000000000000000000000000000000d000a2400000000000000000000000000000000000000000d008f2d00000000000000000000000000000000000000000d002d1100000000000000000000000000000000000000000c00f00f00000000000000000000000000000000000000000c00201000000000000000000000000000000000000000000c00501000000000000000000000000000000000000000000d00f10600000000000000000000000000000000000000000d00033800000000000000000000000000000000000000000d00e12e00000000000000000000000000000000000000000d006a1900000000000000000000000000000000000000000d00731900000000000000000000000000000000000000000d00142f00000000000000000000000000000000000000000d00721600000000000000000000000000000000000000000d00084800000000000000000000000000000000000000000400406e010000000000000000000000000000000000000004004e6e010000000000000000000000000000000000000004002eb30100000000000000000000000000000000000000040030b30100000000000000000000000000000000000000040072b40100000000000000000000000000000000000000040056b601000000000000000000000000000000000000000400acb60100000000000000000000000000000000000000040024ba0100000000000000000000000000000000000000040032ba01000000000000000000000000000000000000000400b0bb01000000000000000000000000000000000000000400c2bb01000000000000000000000000000000000000000400d4bb01000000000000000000000000000000000000000400e2bb01000000000000000000000000000000000000000400f0bb01000000000000000000000000000000000000000400febb010000000000000000000000000000000000000004006ebc010000000000000000000000000000000000000004002abe01000000000000000000000000000000000000000400debe0100000000000000000000000000000000000000040016bf0100000000000000000000000000000000000000040020bf01000000000000000000000000000000000000000400d6bf0100000000000000000000000000000000000000040010c00100000000000000000000000000000000000000040030c10100000000000000000000000000000000000000040030c201000000000000000000000000000000000000000400c8c201000000000000000000000000000000000000000400d6c20100000000000000000000000000000000000000040048c301000000000000000000000000000000000000000400bac301000000000000000000000000000000000000000400d0c30100000000000000000000000000000000000000040072c401000000000000000000000000000000000000000400e2c401000000000000000000000000005a6900000400f1ff00000000000000000000000000000000686900000200040092940200000000003e000000000000006f69000000000400929402000000000000000000000000007269000002000400d0940200000000000e000000000000008569000000000400d0940200000000000000000000000000886900000100070098ca02000000000008000000000000009369000002000400de94020000000000c21a000000000000a469000000000400de940200000000000000000000000000a769000002000400a0af020000000000ae00000000000000bd69000000000400a0af0200000000000000000000000000c0690000000004004eb00200000000000000000000000000c369000000000400f0b00200000000000000000000000000c66900000000040042b10200000000000000000000000000c96900000000040058b10200000000000000000000000000cc69000000000400d2940200000000000000000000000000d1690000000004002c950200000000000000000000000000d66900000000040040950200000000000000000000000000db6900000000040088950200000000000000000000000000e0690000000004009a950200000000000000000000000000e569000000000400ec950200000000000000000000000000ea69000000000400f4950200000000000000000000000000ef6900000000040046960200000000000000000000000000f46900000000040050960200000000000000000000000000f96900000000040004950200000000000000000000000000fd690000000004006caf0200000000000000000000000000016a0000000004000cb00200000000000000000000000000066a00000000040030b002000000000000000000000000000b6a00000000040002b00200000000000000000000000000106a0000000004006cb00200000000000000000000000000156a00000000040076b002000000000000000000000000001a6a00000000040080b002000000000000000000000000001f6a0000000004008ab00200000000000000000000000000246a00000000040094b00200000000000000000000000000296a0000000004009eb002000000000000000000000000002e6a000000000400a8b00200000000000000000000000000336a000000000400b2b00200000000000000000000000000386a000000000400c2b002000000000000000000000000003d6a00000000040034b10200000000000000000000000000426a00000000040054b10200000000000000000000000000476a00000000040024b202000000000000000000000000004c6a000000000400a2b10200000000000000000000000000516a000000000400cab10200000000000000000000000000566a00000400f1ff000000000000000000000000000000005c6a00000000040030b202000000000000000000000000005f6a000000000400feb20200000000000000000000000000626a00000000040026b70200000000000000000000000000656a0000000004004cb70200000000000000000000000000686a000000000400fcb202000000000000000000000000006c6a000000000400ecb20200000000000000000000000000706a00000000040022b70200000000000000000000000000756a000000000400dab302000000000000000000000000007a6a00000000040022b302000000000000000000000000007f6a000000000400c4b50200000000000000000000000000846a0000000004001eb30200000000000000000000000000896a000000000400eeb302000000000000000000000000008e6a0000000004009ab30200000000000000000000000000936a00000000040058b30200000000000000000000000000986a0000000004005cb602000000000000000000000000009d6a00000000040068b30200000000000000000000000000a26a000000000400c0b30200000000000000000000000000a76a000000000400ccb30200000000000000000000000000ac6a000000000400aeb50200000000000000000000000000b16a000000000400a2b40200000000000000000000000000b66a0000000004008cb60200000000000000000000000000bb6a000000000400ceb50200000000000000000000000000c06a00000000040038b40200000000000000000000000000c56a0000000004003cb50200000000000000000000000000ca6a00000000040084b50200000000000000000000000000cf6a000000000400aab50200000000000000000000000000d46a000000000400d0b30200000000000000000000000000d96a000000000400f0b50200000000000000000000000000de6a00000000040066b60200000000000000000000000000e36a000000000400b6b60200000000000000000000000000e86a00000000040036b30200000000000000000000000000ed6a0000000004003cb70200000000000000000000000000f36a00000000040040b70200000000000000000000000000f96a00000000040028b70200000000000000000000000000ff6a0000000004002cb80200000000000000000000000000056b0000000004000cb902000000000000000000000000000b6b00000000040030b80200000000000000000000000000116b00000000040098b80200000000000000000000000000176b00000000040012b902000000000000000000000000001d6b0000000004000eb90200000000000000000000000000236b000000000400aeb70200000000000000000000000000296b00000000040082b802000000000000000000000000002f6b00000000040028b90200000000000000000000000000356b0000000004004eb802000000000000000000000000003b6b00000000040048b80200000000000000000000000000416b00000000040018b90200000000000000000000000000476b0000000004006cb802000000000000000000000000004d6b0000000004002cb90200000000000000000000000000536b000000000400b0b80200000000000000000000000000596b000000000400aab802000000000000000000000000005f6b0000000004001cb90200000000000000000000000000656b000000000400d8b802000000000000000000000000006b6b000000000400fab80200000000000000000000000000716b000000000400f8b80200000000000000000000000000776b000000000400f4b802000000000000000000000000007d6b00000000040062b80200000000000000000000000000836b000000000400c2b802000000000000000000000000009f6b0000020204004cb7020000000000e601000000000000a76b000002020400feb20200000000002804000000000000ae6b00000202040026b70200000000002600000000000000b56b00000202040030b2020000000000ce00000000000000896b000012000400e0470100000000009025000000000000986b00001000040074360100000000000000000000000000bc6b00001200040042b10200000000001600000000000000cb6b00001200040058b1020000000000d800000000000000d96b000012000400f0b00200000000005200000000000000f56b0000120004004eb0020000000000a200000000000000002e726f64617461002e73726f646174612e63737438002e65685f6672616d65002e74657874002e7364617461002e64617461002e73646174612e6d656d7365745f762e30002e627373002e64656275675f616262726576002e64656275675f696e666f002e64656275675f6172616e676573002e64656275675f72616e676573002e64656275675f737472002e64656275675f7075626e616d6573002e64656275675f7075627479706573002e72697363762e61747472696275746573002e64656275675f6c696e65002e636f6d6d656e74002e73796d746162002e7368737472746162002e73747274616200007374616b655f736d742e646436616664343835633633343335632d6367752e30002e4c435049305f30005f5a4e34636f72653370747231373364726f705f696e5f706c616365244c5424616c6c6f632e2e7665632e2e696e746f5f697465722e2e496e746f49746572244c5424244c502424753562247538247533622424753230243230247535642424432424753562247538247533622424753230243332247535642424432461786f6e5f74797065732e2e67656e6572617465642e2e7374616b655f7265616465722e2e5374616b65496e666f44656c74612452502424475424244754243137683236336137653365303866636139333745002e4c706372656c5f686930005f5a4e36345f244c5424616c6c6f632e2e72632e2e5263244c54245424475424247532302461732475323024636f72652e2e6f70732e2e64726f702e2e44726f70244754243464726f703137683663346239333364656266363135663545005f5f727573745f6465616c6c6f63005f5a4e34636f726533707472343664726f705f696e5f706c616365244c5424616c6c6f632e2e7665632e2e566563244c5424753824475424244754243137683361313733353239636533623265663445005f5a4e34636f726533707472383864726f705f696e5f706c616365244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e7365742e2e4254726565536574244c54247574696c2e2e736d742e2e4c6f636b496e666f24475424244754243137683665343465643866393463343166666345002e4c706372656c5f686931002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e30005f5a4e34636f72653970616e69636b696e673570616e69633137686437373538656430613265383739363145005f5a4e35616c6c6f633131636f6c6c656374696f6e733562747265653373657432314254726565536574244c542454244324412447542436696e736572743137686464393035633939376636373034323545005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565367365617263683134325f244c5424696d706c2475323024616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e4e6f6465526566244c5424426f72726f77547970652443244b24432456244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4c6561664f72496e7465726e616c244754242447542431317365617263685f747265653137683334313732383863663534343435313045005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f646532314c6561664e6f6465244c54244b2443245624475424336e65773137683030343135616633666232326365633045005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f64653235496e7465726e616c4e6f6465244c54244b2443245624475424336e65773137683032323863313432336565363266306545005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f646532313448616e646c65244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e4e6f6465526566244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4d75742443244b24432456244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e496e7465726e616c24475424244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e45646765244754243130696e736572745f6669743137686333643836376265346235366332393945002e4c706372656c5f686934002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3639002e4c706372656c5f686935002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3635005f5a4e34636f726535736c69636532395f244c5424696d706c24753230242475356224542475356424244754243135636f70795f66726f6d5f736c69636531376c656e5f6d69736d617463685f6661696c3137686531663934356265353831313135613845002e4c706372656c5f686936002e4c706372656c5f686932002e4c706372656c5f686933002e4c706372656c5f686937002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3537002e4c706372656c5f686938005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f64653132354e6f6465526566244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4d75742443244b24432456244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4c6561664f72496e7465726e616c24475424313663686f6f73655f706172656e745f6b763137683139343665383636343762653264393545005f5a4e34636f72653970616e69636b696e67313870616e69635f6e6f756e77696e645f666d743137683133386130386530383963323036303445005f5f727573745f616c6c6f63005f5f727573745f616c6c6f635f6572726f725f68616e646c6572005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b2443245624475424313562756c6b5f737465616c5f6c6566743137686539616634316334303135636434623645002e4c706372656c5f686939002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3733002e4c706372656c5f68693131002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3735002e4c706372656c5f68693130002e4c706372656c5f68693132002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3737005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b2443245624475424313662756c6b5f737465616c5f72696768743137686162393832373662656263346330393645002e4c706372656c5f68693133002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3830002e4c706372656c5f68693135002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3832002e4c706372656c5f68693134002e4c706372656c5f68693136005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b244324562447542432356d657267655f747261636b696e675f6368696c645f656467653137683538306266633666353961646136383045002e4c706372656c5f68693138002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3835002e4c706372656c5f68693137002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3837005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b244324562447542438646f5f6d657267653137683762346633316135393139303638643245002e4c706372656c5f68693139005f5a4e35616c6c6f633131636f6c6c656374696f6e733562747265653672656d6f76653235395f244c5424696d706c2475323024616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e48616e646c65244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e4e6f6465526566244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4d75742443244b24432456244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4c65616624475424244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4b562447542424475424313472656d6f76655f6c6561665f6b763137683034323333323932386162316238636645002e4c706372656c5f68693230005f5a4e37636b625f73746433656e7634415247563137683036373561626564353032343439613545005f5a4e37636b625f7374643130686967685f6c6576656c31316c6f61645f7363726970743137683962326234613433643962613162666545005f5a4e3131636b625f747970655f696431366861735f747970655f69645f63656c6c3137683163316466616433653431643434383645005f5a4e38345f244c54247574696c2e2e6572726f722e2e4572726f72247532302461732475323024636f72652e2e636f6e766572742e2e46726f6d244c5424636b625f747970655f69642e2e4572726f7224475424244754243466726f6d3137683537363538306531656461613935643645005f5a4e347574696c3668656c706572313663616c635f7363726970745f686173683137686361393462346333346566393134393545005f5a4e35616c6c6f63377261775f7665633139526177566563244c54245424432441244754243131616c6c6f636174655f696e3137683961373435623837316432623838663945005f5a4e347574696c3668656c70657232376765745f63656c6c5f636f756e745f62795f747970655f686173683137683636366663636666636434353161366445005f5a4e37636b625f7374643130686967685f6c6576656c31396c6f61645f63656c6c5f747970655f686173683137686661353738353337303831333261613945005f5a4e39305f244c54247574696c2e2e6572726f722e2e4572726f72247532302461732475323024636f72652e2e636f6e766572742e2e46726f6d244c5424636b625f7374642e2e6572726f722e2e5379734572726f7224475424244754243466726f6d3137686233643163343538633564356263343545002e4c706372656c5f68693234002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e383436002e4c706372656c5f68693236005f5a4e37636b625f7374643130686967685f6c6576656c31306c6f61645f696e7075743137686333316231653162623031363962653245002e4c706372656c5f68693233005f5a4e3130626c616b6532625f727337626c616b6532623134426c616b6532624275696c646572356275696c643137683463643438663738663037316532306145002e4c706372656c5f68693235005f5a4e34636f726533707472353564726f705f696e5f706c616365244c54246d6f6c6563756c652e2e6572726f722e2e566572696669636174696f6e4572726f72244754243137683936383830623737653965663033383845002e4c706372656c5f68693237002e4c706372656c5f68693238002e4c706372656c5f68693239002e4c706372656c5f68693231007374722e342e3733005f5a4e34636f726535736c69636535696e64657837345f244c5424696d706c2475323024636f72652e2e6f70732e2e696e6465782e2e496e646578244c542449244754242475323024666f72247532302424753562245424753564242447542435696e6465783137683064326565363561653136626361336545005f5a4e3131315f244c5424616c6c6f632e2e7665632e2e566563244c54245424475424247532302461732475323024616c6c6f632e2e7665632e2e737065635f66726f6d5f697465725f6e65737465642e2e5370656346726f6d497465724e6573746564244c5424542443244924475424244754243966726f6d5f697465723137683032353562336632346332623633633445005f5a4e35616c6c6f63337665633136566563244c542454244324412447542434707573683137683832346530366138613965323339383745005f5a4e34636f7265346974657236747261697473386974657261746f72384974657261746f7233616e793137683031323866356465313834336464653445002e4c706372656c5f68693331002e4c706372656c5f68693232007374722e302e313130002e4c706372656c5f68693330005f5a4e3130325f244c5424636b625f7374616e64616c6f6e655f74797065732e2e67656e6572617465642e2e626c6f636b636861696e2e2e42797465735265616465722475323024617324753230246d6f6c6563756c652e2e7072656c7564652e2e52656164657224475424367665726966793137683135663233383466353032373265326345005f5a4e386d6f6c6563756c6535627974657335427974657335736c6963653137683133633337653065643765643238336345005f5a4e3230636b625f7374616e64616c6f6e655f74797065733967656e6572617465643130626c6f636b636861696e354279746573387261775f646174613137686165613062386538653731396665363945005f5a4e347574696c3668656c70657231386765745f7374616b655f736d745f646174613137683531393538393938623361383432363145005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231365374616b65536d7443656c6c4461746131366d657461646174615f747970655f69643137683333316537333761333766666465306145005f5a4e347574696c3668656c70657231326765745f747970655f6964733137683161323938396534376363663639393545005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f72656164657237547970654964733134787564745f747970655f686173683137686334653636633566343738343237356145005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f726561646572375479706549647331397374616b655f736d745f636f64655f686173683137683939313230643232643561376161363745005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f726561646572375479706549647331377374616b655f736d745f747970655f69643137683133613730383736373561386135323245005f5a4e347574696c3668656c70657231356765745f7363726970745f686173683137683861333134336361336163636135633445005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f72656164657237547970654964733230636865636b706f696e745f636f64655f686173683137683561366363373337366465333564383045005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f72656164657237547970654964733138636865636b706f696e745f747970655f69643137683062376537323033303666383865346345005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f7265616465723754797065496473313877697468647261775f636f64655f686173683137686636356461336666633664366137323445005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f726561646572375479706549647331386d657461646174615f636f64655f686173683137683263623137613437626166656264306645005f5a4e313061786f6e5f74797065733967656e65726174656431356d657461646174615f726561646572375479706549647331366d657461646174615f747970655f69643137683833306539326563613930383864363745005f5a4e3230636b625f7374616e64616c6f6e655f74797065733967656e6572617465643130626c6f636b636861696e31315769746e65737341726773346c6f636b3137686233326333343036613431316531636245005f5a4e39385f244c54246d6f6c6563756c65322e2e7265616465722e2e437572736f72247532302461732475323024636f72652e2e636f6e766572742e2e46726f6d244c5424616c6c6f632e2e7665632e2e566563244c542475382447542424475424244754243466726f6d3137686365383937663564613837343036643045005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231345374616b65496e666f44656c7461313169735f696e6372656173653137683166386136356661303836623163316645005f5a4e347574696c3668656c70657231376765745f63757272656e745f65706f63683137683433313039626562306665666534313945005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231385374616b65536d74557064617465496e666f3135616c6c5f7374616b655f696e666f733137686331656532343334363962343463366245005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231305374616b65496e666f73336c656e3137683862303137666338646362303233393945005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231305374616b65496e666f73336765743137683536663765343736643831623335613045005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f726561646572395374616b65496e666f34616464723137683737663935343236353164653934373045005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231345374616b65496e666f44656c746136616d6f756e743137683736303137613463316430633135626445005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231385374616b65536d74557064617465496e666f31356f6c645f65706f63685f70726f6f663137683835396638343561623737663561346545005f5a4e347574696c33736d7431317536345f746f5f683235363137683630616266646338653134653935363145005f5a4e347574696c33736d7431377665726966795f326c617965725f736d743137683133343062636139316137313632616545005f5a4e347574696c3668656c70657232326765745f7374616b655f7570646174655f696e666f733137686337343437303336323761616365383045005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231345374616b65496e666f44656c74613138696e61756775726174696f6e5f65706f63683137683538323561303933383837366165313345005f5a4e347574696c3668656c70657233306765745f7374616b655f61745f646174615f62795f6c6f636b5f686173683137683536356232313136353933333665623945005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231355374616b65417443656c6c446174613564656c74613137683762333332613765343438316530613845005f5a4e3130385f244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6d61702e2e49746572244c54244b2443245624475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683932393561376437613164316266393145005f5a4e347574696c3668656c706572323563616c635f7769746864726177616c5f6c6f636b5f686173683137683038613966633761623133353165326345005f5a4e347574696c3668656c70657233336765745f77697468647261775f61745f646174615f62795f6c6f636b5f686173683137686531356438613763623138663661663445005f5a4e347574696c3668656c70657231356765745f71756f72756d5f73697a653137683930353932376137656234333038306645005f5a4e313061786f6e5f74797065733967656e65726174656431327374616b655f72656164657231385374616b65536d74557064617465496e666f31356e65775f65706f63685f70726f6f663137686236623761343265306435646564653745002e4c706372656c5f68693332002e4c706372656c5f68693433007374722e31002e4c706372656c5f68693333002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3436002e4c706372656c5f68693334002e4c616e6f6e2e36633237623166666234666234346562313164656530663863336331326232322e33005f5a4e34636f726536726573756c743133756e777261705f6661696c65643137683030653934303161326339653536633045002e4c706372656c5f68693435002e4c706372656c5f68693436002e4c706372656c5f68693335002e4c706372656c5f68693336002e4c616e6f6e2e36633237623166666234666234346562313164656530663863336331326232322e32002e4c706372656c5f68693337002e4c706372656c5f68693338002e4c706372656c5f68693339002e4c706372656c5f68693430002e4c706372656c5f68693431002e4c706372656c5f68693432002e4c706372656c5f68693434002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e363300727573745f626567696e5f756e77696e64005f5a4e37636b625f7374643873797363616c6c73366e617469766534657869743137683163616638653234666532613530323145005f5f72675f616c6c6f63005f5a4e3130365f244c542462756464795f616c6c6f632e2e6e6f6e5f746872656164736166655f616c6c6f632e2e4e6f6e54687265616473616665416c6c6f63247532302461732475323024636f72652e2e616c6c6f632e2e676c6f62616c2e2e476c6f62616c416c6c6f632447542435616c6c6f633137683966656332343337626566343266383945005f5f72675f6465616c6c6f63005f5a4e3130365f244c542462756464795f616c6c6f632e2e6e6f6e5f746872656164736166655f616c6c6f632e2e4e6f6e54687265616473616665416c6c6f63247532302461732475323024636f72652e2e616c6c6f632e2e676c6f62616c2e2e476c6f62616c416c6c6f6324475424376465616c6c6f633137686530336235656339643238613732396445005f5f72675f7265616c6c6f63005f5f72675f616c6c6f635f7a65726f6564005f5f727573745f7265616c6c6f63005f5f727573745f616c6c6f635f7a65726f6564005f5f72646c5f6f6f6d005f5a4e35616c6c6f63377261775f766563313763617061636974795f6f766572666c6f773137683736396433373734353939336431626545005f5a4e396d6f6c6563756c65323672656164657236437572736f72323164796e7665635f736c6963655f62795f696e6465783137683464633230383535323662653634303045005f5a4e396d6f6c6563756c6532367265616465723130385f244c5424696d706c2475323024636f72652e2e636f6e766572742e2e46726f6d244c54246d6f6c6563756c65322e2e7265616465722e2e437572736f72244754242475323024666f722475323024616c6c6f632e2e7665632e2e566563244c5424753824475424244754243466726f6d3137683965653331373661666261663535343545002e4c706372656c5f68693437002e4c706372656c5f68693438002e4c616e6f6e2e65383134633736363361666663333138633766356639363865643531663662352e3139002e4c706372656c5f68693439002e4c706372656c5f68693530002e4c706372656c5f68693531002e4c706372656c5f68693532002e4c706372656c5f68693533002e4c706372656c5f68693534002e4c706372656c5f68693535002e4c706372656c5f68693536002e4c706372656c5f68693537002e4c706372656c5f68693538002e4c706372656c5f68693539002e4c706372656c5f68693630002e4c706372656c5f68693631002e4c706372656c5f68693632005f5a4e396d6f6c6563756c65323672656164657238355f244c5424696d706c2475323024636f72652e2e636f6e766572742e2e46726f6d244c54246d6f6c6563756c65322e2e7265616465722e2e437572736f72244754242475323024666f7224753230247538244754243466726f6d3137686461653235633931336631613435396545002e4c706372656c5f68693633002e4c706372656c5f68693634002e4c706372656c5f68693635002e4c706372656c5f68693636005f5a4e396d6f6c6563756c65323672656164657238365f244c5424696d706c2475323024636f72652e2e636f6e766572742e2e46726f6d244c54246d6f6c6563756c65322e2e7265616465722e2e437572736f72244754242475323024666f722475323024753634244754243466726f6d3137686232663035653938653831303635333145002e4c706372656c5f68693637002e4c706372656c5f68693638002e4c706372656c5f68693639002e4c706372656c5f68693730002e4c706372656c5f68693731002e4c706372656c5f68693732002e4c706372656c5f68693733002e4c706372656c5f68693734005f5a4e396d6f6c6563756c65323672656164657236437572736f723876616c69646174653137683930306131623931383065653939313845005f5a4e396d6f6c6563756c65323672656164657236437572736f7231346765745f6974656d5f636f756e743137683362393033346337303939633162346445002e4c706372656c5f68693735002e4c706372656c5f68693736002e4c706372656c5f68693737002e4c706372656c5f68693738002e4c706372656c5f68693739002e4c706372656c5f68693830005f5a4e396d6f6c6563756c65323672656164657236437572736f723139636f6e766572745f746f5f72617762797465733137683634326263616436376665326537643145002e4c706372656c5f68693831002e4c706372656c5f68693832002e4c706372656c5f68693833002e4c706372656c5f68693834002e4c706372656c5f68693835002e4c706372656c5f68693836002e4c706372656c5f68693837002e4c706372656c5f68693838005f5a4e3131626c616b6532625f72656637777261707065723134426c616b6532624275696c646572356275696c643137683964636431366662373535323133626345005f5a4e3131626c616b6532625f7265663131626c616b6532625f7265663138626c616b6532625f696e69745f706172616d3137683431613831343963666239633164343445005f5a4e3131626c616b6532625f7265663131626c616b6532625f7265663134626c616b6532625f7570646174653137683337646637643338333264666265336545002e4c706372656c5f68693839005f5a4e3131626c616b6532625f7265663131626c616b6532625f7265663130626c616b6532625f49563137686532356438333932346363316638393145005f5a4e3131626c616b6532625f7265663131626c616b6532625f7265663136626c616b6532625f636f6d70726573733137683531363361326435303733336262323945002e4c43504934395f30002e4c43504934395f31002e4c43504934395f32002e4c43504934395f33002e4c43504934395f34002e4c43504934395f35002e4c43504934395f36002e4c43504934395f37002e4c706372656c5f68693930002e4c706372656c5f68693931002e4c706372656c5f68693932002e4c706372656c5f68693933002e4c706372656c5f68693934002e4c706372656c5f68693935002e4c706372656c5f68693936002e4c706372656c5f68693937005f5a4e3131626c616b6532625f726566377772617070657237426c616b6532623866696e616c697a653137683431356365303263316365386263623745005f5a4e313162756464795f616c6c6f63313162756464795f616c6c6f6331304275646479416c6c6f63336e65773137683039343964346234353436656265666245005f5a4e313162756464795f616c6c6f63313162756464795f616c6c6f6337726f756e6475703137686533656266373734346663663366363345002e4c706372656c5f6869313035007374722e342e3633005f5a4e313162756464795f616c6c6f63313162756464795f616c6c6f63366e626c6f636b3137683537623963376462363561386133343745005f5a4e313162756464795f616c6c6f63313162756464795f616c6c6f6331304275646479416c6c6f633131626c6f636b5f696e6465783137683333633165376336333564613363643945005f5a4e34636f7265366f7074696f6e31336578706563745f6661696c65643137686332333330616533386638616564396545002e4c706372656c5f6869313130002e4c706372656c5f6869313036002e4c706372656c5f6869313037002e4c706372656c5f68693938002e4c706372656c5f6869313030007374722e322e3634002e4c706372656c5f6869313031007374722e332e3635002e4c706372656c5f6869313032002e4c706372656c5f6869313033007374722e312e3632002e4c706372656c5f6869313034002e4c706372656c5f6869313131002e4c706372656c5f6869313038007374722e302e3631002e4c706372656c5f68693939002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3135002e4c706372656c5f6869313132002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3238005f5a4e34636f72653970616e69636b696e67313370616e69635f646973706c61793137683538303536323433613031393534316645002e4c706372656c5f6869313039002e4c706372656c5f6869313133002e4c706372656c5f6869313134002e4c706372656c5f6869313135002e4c706372656c5f6869313136002e4c706372656c5f6869313137002e4c706372656c5f6869313139002e4c706372656c5f6869313230002e4c706372656c5f6869313138002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3338005f5a4e313162756464795f616c6c6f633130666173745f616c6c6f633946617374416c6c6f63336e65773137683239303962396561363461333531383845002e4c706372656c5f6869313232002e4c706372656c5f6869313231002e4c706372656c5f6869313233002e4c706372656c5f6869313234005f5a4e397374616b655f736d7435414c4c4f433137683263336231343434623861633161633845002e4c706372656c5f6869313238002e4c706372656c5f6869313333002e4c706372656c5f6869313334002e4c706372656c5f6869313331002e4c706372656c5f6869313335002e4c706372656c5f6869313336002e4c706372656c5f6869313332002e4c706372656c5f6869313237002e4c706372656c5f6869313239002e4c706372656c5f6869313330002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e32002e4c706372656c5f6869313235002e4c706372656c5f6869313236002e4c706372656c5f6869313337002e4c706372656c5f6869313338002e4c706372656c5f6869313339002e4c706372656c5f6869313433002e4c706372656c5f6869313432002e4c706372656c5f6869313436002e4c706372656c5f6869313438002e4c706372656c5f6869313439002e4c706372656c5f6869313530002e4c706372656c5f6869313437002e4c706372656c5f6869313430002e4c706372656c5f6869313431002e4c706372656c5f6869313434002e4c706372656c5f6869313435005f5a4e35616c6c6f63377261775f7665633139526177566563244c54245424432441244754243131616c6c6f636174655f696e3137683334393639363464643031633234363645005f5a4e35616c6c6f63377261775f7665633139526177566563244c542454244324412447542437726573657276653231646f5f726573657276655f616e645f68616e646c653137686234636364626536643135363830353445002e4c706372656c5f6869313531007374722e302e3731005f5a4e35616c6c6f63377261775f7665633139526177566563244c5424542443244124475424313467726f775f616d6f7274697a65643137683131313435313531653037646531613245005f5a4e35616c6c6f63377261775f766563313166696e6973685f67726f773137683362363537323731663362336132663345005f5a4e35616c6c6f63377261775f7665633139526177566563244c54245424432441244754243136726573657276655f666f725f707573683137683364383734353931323332303230376445002e4c706372656c5f6869313532002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e313734002e4c706372656c5f6869313533002e4c706372656c5f6869313534005f5a4e3230636b625f7374616e64616c6f6e655f74797065733130636f6e76657273696f6e3130626c6f636b636861696e3134395f244c5424696d706c2475323024636b625f7374616e64616c6f6e655f74797065732e2e7072656c7564652e2e5061636b244c5424636b625f7374616e64616c6f6e655f74797065732e2e67656e6572617465642e2e626c6f636b636861696e2e2e427974653332244754242475323024666f72247532302424753562247538247533622424753230243332247535642424475424347061636b3137683838633365666265633136666335636345005f5a4e3230636b625f7374616e64616c6f6e655f74797065733130636f6e76657273696f6e397072696d69746976653133365f244c5424696d706c2475323024636b625f7374616e64616c6f6e655f74797065732e2e7072656c7564652e2e5061636b244c5424636b625f7374616e64616c6f6e655f74797065732e2e67656e6572617465642e2e626c6f636b636861696e2e2e4279746573244754242475323024666f72247532302424753562247538247535642424475424347061636b3137686534363231633861323935306563356145005f5a4e3133325f244c5424616c6c6f632e2e7665632e2e566563244c5424542443244124475424247532302461732475323024616c6c6f632e2e7665632e2e737065635f657874656e642e2e53706563457874656e64244c54242452462454244324636f72652e2e736c6963652e2e697465722e2e49746572244c5424542447542424475424244754243131737065635f657874656e643137683464663561353366366631653763336445002e4c706372656c5f6869313535007374722e322e3730005f5a4e39375f244c5424636b625f7374616e64616c6f6e655f74797065732e2e67656e6572617465642e2e626c6f636b636861696e2e2e5363726970742475323024617324753230246d6f6c6563756c652e2e7072656c7564652e2e456e746974792447542431316e65775f6275696c6465723137683663323863633439326130386634363645005f5a4e3130355f244c5424636b625f7374616e64616c6f6e655f74797065732e2e67656e6572617465642e2e626c6f636b636861696e2e2e5363726970744275696c6465722475323024617324753230246d6f6c6563756c652e2e7072656c7564652e2e4275696c64657224475424356275696c643137683462313334356436646334623638326145002e4c706372656c5f6869313536002e4c706372656c5f6869313537002e4c706372656c5f6869313538005f5a4e36315f244c5424636b625f7374642e2e6572726f722e2e5379734572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683863383033303266623836336136303845002e4c706372656c5f6869313539002e4c4a544937365f30002e4c424237365f31002e4c706372656c5f6869313630002e4c616e6f6e2e34313466363731613135666237623063306532636261396133343630323939342e3339002e4c424237365f32002e4c706372656c5f6869313631002e4c616e6f6e2e34313466363731613135666237623063306532636261396133343630323939342e3338002e4c424237365f33002e4c706372656c5f6869313632002e4c616e6f6e2e34313466363731613135666237623063306532636261396133343630323939342e3336002e4c706372656c5f6869313633002e4c616e6f6e2e34313466363731613135666237623063306532636261396133343630323939342e3337002e4c424237365f34002e4c706372656c5f6869313634002e4c424237365f36002e4c706372656c5f6869313635002e4c616e6f6e2e34313466363731613135666237623063306532636261396133343630323939342e3333002e4c706372656c5f6869313636002e4c616e6f6e2e34313466363731613135666237623063306532636261396133343630323939342e3334005f5a4e34636f726533666d7439466f726d6174746572323564656275675f7475706c655f6669656c64315f66696e6973683137683963326264643732306464613133376545005f5a4e34636f726533707472323864726f705f696e5f706c616365244c542424524624753634244754243137683536663832373834643464373061633345002e4c706372656c5f6869313637002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e343734005f5a4e37636b625f7374643130686967685f6c6576656c31396c6f61645f63656c6c5f6c6f636b5f686173683137686238376330343133623735373432633545005f5a4e37636b625f7374643130686967685f6c6576656c31346c6f61645f63656c6c5f646174613137686438663961623933373437336639633645002e4c706372656c5f6869313638002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e343330002e4c706372656c5f6869313730002e4c706372656c5f6869313639002e4c706372656c5f6869313731002e4c706372656c5f6869313732002e4c706372656c5f6869313733002e4c706372656c5f6869313735002e4c706372656c5f6869313734002e4c706372656c5f6869313736002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e3936002e4c706372656c5f6869313737002e4c616e6f6e2e65653231316338393139316237376236333039663861393366623935653339352e3234005f5a4e34636f7265336f70733866756e6374696f6e36466e4f6e63653963616c6c5f6f6e63653137683331326365396462383432326365623645005f5a4e34636f72653370747231303264726f705f696e5f706c616365244c542424524624636f72652e2e697465722e2e61646170746572732e2e636f706965642e2e436f70696564244c5424636f72652e2e736c6963652e2e697465722e2e49746572244c542475382447542424475424244754243137683465633534623435323134663763393045002e4c43504938385f30005f5a4e34636f726533666d74336e756d33696d7037666d745f7536343137683238366534643532373433386334363745002e4c706372656c5f6869313738002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333234002e4c706372656c5f6869313739002e4c706372656c5f6869313830002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3233005f5a4e34636f726533666d7439466f726d617474657231327061645f696e74656772616c3137686238656639343965396131613633346545005f5a4e34636f726533666d7439466f726d617474657231327061645f696e74656772616c313277726974655f7072656669783137683834663538656430383761336264393345002e4c43504939315f30002e4c43504939315f31005f5a4e34636f726533666d7439466f726d6174746572337061643137683433336537613934646232626438653245002e4c706372656c5f6869313831002e4c706372656c5f6869313832005f5a4e34636f726533666d743577726974653137683537653362636463656237646630393145002e4c706372656c5f6869313833005f5a4e36305f244c5424636f72652e2e63656c6c2e2e426f72726f774572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137686163386261333334363731373261333845002e4c706372656c5f6869313834002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e313730005f5a4e36335f244c5424636f72652e2e63656c6c2e2e426f72726f774d75744572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683636336332373865383138373636393045002e4c706372656c5f6869313835002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e313731005f5a4e34636f726533666d74336e756d35335f244c5424696d706c2475323024636f72652e2e666d742e2e4c6f7765724865782475323024666f7224753230246936342447542433666d743137686632356530653835343735353364373145002e4c706372656c5f6869313836002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333232002e4c4350493130305f30002e4c4350493130305f31002e4c4350493130305f32005f5a4e36385f244c5424636f72652e2e666d742e2e6275696c646572732e2e50616441646170746572247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f7374723137686539366438303337316562386433343445002e4c706372656c5f6869313837002e4c706372656c5f6869313838002e4c706372656c5f6869313839002e4c706372656c5f6869313930005f5a4e34636f726533666d74355772697465313077726974655f636861723137686664666234386663643336373461323845005f5a4e34636f726533666d743557726974653977726974655f666d743137683364623431343565346436363932376245002e4c706372656c5f6869313931002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333237005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f7374723137683865303931326361326264646233386345005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e577269746524475424313077726974655f636861723137683239666437616639333939643762333645005f5a4e35305f244c5424245246246d7574247532302457247532302461732475323024636f72652e2e666d742e2e5772697465244754243977726974655f666d743137683565373464633863623261616161323645002e4c706372656c5f6869313932005f5a4e34636f726533666d74386275696c64657273313044656275675475706c65356669656c643137686134393061356537663734366534656245002e4c706372656c5f6869313934002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e323933002e4c706372656c5f6869313935002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333030002e4c706372656c5f6869313933002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333031002e4c706372656c5f6869313936002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e323839002e4c706372656c5f6869313937002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e323932005f5a4e34636f726533666d74386275696c6465727338446562756753657435656e7472793137686531623638303262326163636539656445002e4c706372656c5f6869323031002e4c706372656c5f6869313939002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333033002e4c706372656c5f6869313938002e4c706372656c5f6869323030002e4c706372656c5f6869323033002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333032002e4c706372656c5f6869323032002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e313537005f5a4e34636f726533666d74336e756d35325f244c5424696d706c2475323024636f72652e2e666d742e2e55707065724865782475323024666f72247532302469382447542433666d743137683438643832613435336137306166353745002e4c706372656c5f6869323034005f5a4e34636f726533666d74336e756d35325f244c5424696d706c2475323024636f72652e2e666d742e2e4c6f7765724865782475323024666f72247532302469382447542433666d743137683039663834613031663936303437366145002e4c706372656c5f6869323035005f5a4e34325f244c54242452462454247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137686332303631326561373836393861653445002e4c706372656c5f6869323036002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333337005f5a4e36375f244c5424636f72652e2e61727261792e2e54727946726f6d536c6963654572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683532646436363362353834636335356645002e4c706372656c5f6869323037002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e353537002e4c706372656c5f6869323038002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e353333002e4c706372656c5f6869323130002e4c706372656c5f6869323039005f5a4e34636f726533666d74336e756d35335f244c5424696d706c2475323024636f72652e2e666d742e2e55707065724865782475323024666f7224753230246936342447542433666d743137683464336136353331313038303933376445002e4c706372656c5f6869323131005f5a4e35616c6c6f63377261775f7665633139526177566563244c542454244324412447542437726573657276653231646f5f726573657276655f616e645f68616e646c653137686332663335393562613638613033633645005f5a4e34325f244c54242452462454247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683035646461313430303562373034353645005f5a4e34325f244c54242452462454247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683431323134373832613466363464656645005f5a4e36355f244c5424616c6c6f632e2e7665632e2e566563244c5424542443244124475424247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137686464613861616433336135376363313045002e4c706372656c5f6869323132002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e323533002e4c706372656c5f6869323133002e4c706372656c5f6869323134002e4c616e6f6e2e39616236623536633861336165336331383834656237326561613362336632392e333038005f5a4e35616c6c6f63337665633136566563244c54245424432441244754243131657874656e645f776974683137683935323361376565386561616133316645005f5a4e35616c6c6f63377261775f7665633139526177566563244c542454244324412447542437726573657276653231646f5f726573657276655f616e645f68616e646c653137686534386235666233366361343936633545005f5a4e35616c6c6f63377261775f766563313166696e6973685f67726f773137686465323762646133633136313431313345005f5a4e396d6f6c6563756c65323672656164657237726561645f61743137686436323832346538376630396538383045002e4c706372656c5f6869323234007374722e312e333135002e4c706372656c5f6869323137002e4c706372656c5f6869323138002e4c706372656c5f6869323135002e4c706372656c5f6869323136002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e31002e4c706372656c5f6869323233002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3136002e4c706372656c5f6869323235002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3139002e4c706372656c5f6869323139002e4c706372656c5f6869323230002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e36002e4c706372656c5f6869323231002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3132002e4c706372656c5f6869323232002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3134005f5a4e36315f244c54246d6f6c6563756c65322e2e7265616465722e2e4572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683238346238363235356264316239336545002e4c706372656c5f6869323236002e4c7377697463682e7461626c652e5f5a4e36315f244c54246d6f6c6563756c65322e2e7265616465722e2e4572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d743137683238346238363235356264316239336545002e4c706372656c5f6869323237002e4c7377697463682e7461626c652e5f5a4e36315f244c54246d6f6c6563756c65322e2e7265616465722e2e4572726f72247532302461732475323024636f72652e2e666d742e2e44656275672447542433666d7431376832383462383632353562643162393365452e343330002e4c706372656c5f6869323330002e4c706372656c5f6869323238002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e32002e4c706372656c5f6869323239002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e33002e4c706372656c5f6869323331002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3238005f5a4e396d6f6c6563756c65323672656164657236437572736f723133756e7061636b5f6e756d6265723137683635326430373132666263326536343145002e4c706372656c5f6869323332002e4c706372656c5f6869323333002e4c706372656c5f6869323334002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3331002e4c706372656c5f6869323335002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3335002e4c706372656c5f6869323432002e4c706372656c5f6869323336002e4c706372656c5f6869323337002e4c706372656c5f6869323431002e4c706372656c5f6869323338002e4c706372656c5f6869323339002e4c706372656c5f6869323430002e4c706372656c5f6869323433002e4c706372656c5f6869323434002e4c706372656c5f6869323435002e4c706372656c5f6869323436002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3430002e4c706372656c5f6869323437002e4c706372656c5f6869323438002e4c706372656c5f6869323439002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3538002e4c706372656c5f6869323530002e4c706372656c5f6869323531002e4c706372656c5f6869323532002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3634005f5a4e36395f244c5424616c6c6f632e2e7665632e2e566563244c54247538244754242475323024617324753230246d6f6c6563756c65322e2e7265616465722e2e526561642447542434726561643137683538323363346134366134643066373445002e4c706372656c5f6869323533002e4c706372656c5f6869323534002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3638005f5a4e34636f726533707472343664726f705f696e5f706c616365244c5424616c6c6f632e2e7665632e2e566563244c5424753824475424244754243137683139303635656264313265376238616645005f5a4e31387370617273655f6d65726b6c655f74726565346832353634483235363131706172656e745f706174683137683635373836666235326663646564306445005f5a4e37305f244c54247370617273655f6d65726b6c655f747265652e2e747265652e2e4272616e63684b6579247532302461732475323024636f72652e2e636d702e2e4f72642447542433636d703137683263653439633663323334323262346545005f5a4e39385f244c5424636b625f7374642e2e686967685f6c6576656c2e2e517565727949746572244c54244624475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137686231366136333531633137303061613745002e4c706372656c5f6869323535007374722e302e333530002e4c706372656c5f6869323537002e4c706372656c5f6869323536005f5a4e35616c6c6f6335626f7865643136426f78244c542454244324412447542431336e65775f756e696e69745f696e3137683834373362316265336534316438633545005f5a4e35616c6c6f6335626f7865643136426f78244c542454244324412447542431336e65775f756e696e69745f696e3137683761393538346163663734633633393245005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f646532313448616e646c65244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e4e6f6465526566244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4d75742443244b24432456244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e496e7465726e616c24475424244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e45646765244754243130696e736572745f6669743137686530613963663030393033343261333745005f5a4e35616c6c6f633131636f6c6c656374696f6e733562747265653673656172636839315f244c5424696d706c2475323024616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e4e6f6465526566244c5424426f72726f77547970652443244b24432456244324547970652447542424475424313466696e645f6b65795f696e6465783137683538623066623732343130626338653045005f5a4e35616c6c6f633131636f6c6c656374696f6e733562747265653672656d6f76653235395f244c5424696d706c2475323024616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e48616e646c65244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e4e6f6465526566244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4d75742443244b24432456244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4c65616624475424244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4b562447542424475424313472656d6f76655f6c6561665f6b763137683932356266653833663964336631323045005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b244324562447542432356d657267655f747261636b696e675f6368696c645f656467653137683565316662626261313330613939366445005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b2443245624475424313662756c6b5f737465616c5f72696768743137683134353762643930393139373763616445005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b2443245624475424313562756c6b5f737465616c5f6c6566743137686637323766663464373765333137663345005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b244324562447542438646f5f6d657267653137683764663761343032346566636539366545002e4c706372656c5f6869323538002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3731002e4c706372656c5f6869323539002e4c706372656c5f6869323631002e4c706372656c5f6869323630002e4c706372656c5f6869323632002e4c706372656c5f6869323634002e4c706372656c5f6869323633002e4c706372656c5f6869323635002e4c706372656c5f6869323636002e4c706372656c5f6869323638002e4c706372656c5f6869323637002e4c706372656c5f6869323639002e4c706372656c5f6869323730005f5a4e35616c6c6f6335626f7865643136426f78244c542454244324412447542431336e65775f756e696e69745f696e3137683865303536326639626532336432623745005f5a4e35616c6c6f6335626f7865643136426f78244c542454244324412447542431336e65775f756e696e69745f696e3137686630333839343435343838663831633145005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f646532313448616e646c65244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e4e6f6465526566244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4d75742443244b24432456244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e496e7465726e616c24475424244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e45646765244754243130696e736572745f6669743137683463363562306630323863663661333845005f5a4e35616c6c6f633131636f6c6c656374696f6e733562747265653673656172636839315f244c5424696d706c2475323024616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e4e6f6465526566244c5424426f72726f77547970652443244b24432456244324547970652447542424475424313466696e645f6b65795f696e6465783137686366633034636463626438393439336245005f5a4e35616c6c6f633131636f6c6c656374696f6e733562747265653672656d6f76653235395f244c5424696d706c2475323024616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e48616e646c65244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e4e6f6465526566244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4d75742443244b24432456244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4c65616624475424244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4b562447542424475424313472656d6f76655f6c6561665f6b763137686430343065343765356162316639336445005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f64653132354e6f6465526566244c5424616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4d75742443244b24432456244324616c6c6f632e2e636f6c6c656374696f6e732e2e62747265652e2e6e6f64652e2e6d61726b65722e2e4c6561664f72496e7465726e616c24475424313663686f6f73655f706172656e745f6b763137683662323932356361633530363230653245005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b244324562447542432356d657267655f747261636b696e675f6368696c645f656467653137683639343536653266653337656664353245005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b2443245624475424313662756c6b5f737465616c5f72696768743137683333636262626135643162656234643245005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b2443245624475424313562756c6b5f737465616c5f6c6566743137683565653138306237396130613266636245005f5a4e35616c6c6f633131636f6c6c656374696f6e73356274726565346e6f6465323942616c616e63696e67436f6e74657874244c54244b244324562447542438646f5f6d657267653137683062356263386231666365346431343845002e4c706372656c5f6869323731002e4c706372656c5f6869323732002e4c706372656c5f6869323734002e4c706372656c5f6869323733002e4c706372656c5f6869323735002e4c706372656c5f6869323737002e4c706372656c5f6869323736002e4c706372656c5f6869323738002e4c706372656c5f6869323739002e4c706372656c5f6869323831002e4c706372656c5f6869323830002e4c706372656c5f6869323832002e4c706372656c5f6869323833005f5a4e34636f726535736c69636534736f727437726563757273653137686635623239333039636436333933336245005f5a4e34636f726535736c69636534736f72743235696e73657274696f6e5f736f72745f73686966745f6c6566743137683133346537316232363032303439623045005f5a4e34636f726535736c69636534736f72743134627265616b5f7061747465726e733137683038373030316334666161636539623445005f5a4e34636f726535736c69636534736f727432327061727469616c5f696e73657274696f6e5f736f72743137683664666664346137303338356239303045005f5a4e34636f726535736c69636534736f72743868656170736f72743137683739313663343261326535636431383945002e4c4350493136335f30005f5a4e35616c6c6f63377261775f7665633139526177566563244c54245424432441244754243136726573657276655f666f725f707573683137683266373139353338366332346364373445002e4c706372656c5f6869323834005f5a4e31387370617273655f6d65726b6c655f74726565356d65726765356d657267653137683733636631633763646362636630363645002e4c706372656c5f6869323837005f5a4e347574696c33736d7431316e65775f626c616b6532623137686530346638633332383130656566666645005f5a4e31387370617273655f6d65726b6c655f74726565356d6572676531304d6572676556616c756534686173683137686361663934316539633361336137646145002e4c706372656c5f6869323835002e4c706372656c5f6869323836005f5a4e31387370617273655f6d65726b6c655f74726565356d6572676531356d657267655f776974685f7a65726f3137686262316663663731613061663431616545002e4c706372656c5f6869323838002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3331002e4c4350493136395f30002e4c4350493136395f31002e4c4350493136395f32002e4c4350493136395f33002e4c706372656c5f6869323839002e4c706372656c5f6869323930002e4c706372656c5f6869323931002e4c706372656c5f6869323932002e4c706372656c5f6869323933005f5a4e34636f726535736c69636534736f72743236696e73657274696f6e5f736f72745f73686966745f72696768743137686537623533613633393836633665636245002e4c706372656c5f6869323934002e4c4350493137335f30005f5a4e35616c6c6f63377261775f7665633139526177566563244c54245424432441244754243136726573657276655f666f725f707573683137686331393061356231623136306436373545002e4c706372656c5f6869323935005f5a4e39385f244c5424636b625f7374642e2e686967685f6c6576656c2e2e517565727949746572244c54244624475424247532302461732475323024636f72652e2e697465722e2e7472616974732e2e6974657261746f722e2e4974657261746f7224475424346e6578743137683639396362383835316633373032373345002e4c706372656c5f6869323936002e4c706372656c5f6869323937002e4c4a54493137355f30002e4c42423137355f31002e4c42423137355f32002e4c42423137355f33002e4c42423137355f34002e4c42423137355f35002e4c706372656c5f6869323938005f5a4e34636f726533707472373964726f705f696e5f706c616365244c5424636b625f7374616e64616c6f6e655f74797065732e2e67656e6572617465642e2e626c6f636b636861696e2e2e5363726970744275696c646572244754243137683230353465616461363664306463376345002e4c706372656c5f6869323939002e4c706372656c5f6869333030002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3437002e4c706372656c5f6869333032002e4c706372656c5f6869333031002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e313134002e4c706372656c5f6869333033002e4c706372656c5f6869333034002e4c706372656c5f6869333038002e4c706372656c5f6869333035002e4c706372656c5f6869333036002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3438002e4c706372656c5f6869333037002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e313139002e4c706372656c5f6869333132002e4c706372656c5f6869333039002e4c706372656c5f6869333130002e4c706372656c5f6869333131002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e313237002e4c706372656c5f6869333231002e4c706372656c5f6869333133002e4c706372656c5f6869333134002e4c706372656c5f6869333135002e4c706372656c5f6869333136002e4c706372656c5f6869333137002e4c706372656c5f6869333138002e4c706372656c5f6869333139002e4c706372656c5f6869333230002e4c706372656c5f6869333232005f5a4e347574696c3668656c70657232366765745f6d65746164615f646174615f62795f747970655f69643137683437383266333330623964363130353445002e4c706372656c5f6869333235002e4c706372656c5f6869333233002e4c706372656c5f6869333234002e4c706372656c5f6869333236002e4c706372656c5f6869333237002e4c706372656c5f6869333238002e4c706372656c5f6869333239002e4c706372656c5f6869333330002e4c706372656c5f6869333331002e4c706372656c5f6869333332002e4c706372656c5f6869333333002e4c706372656c5f6869333334002e4c706372656c5f6869333335002e4c706372656c5f6869333336002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3532002e4c706372656c5f6869333339002e4c706372656c5f6869333337002e4c706372656c5f6869333338002e4c706372656c5f6869333430002e4c706372656c5f6869333434002e4c706372656c5f6869333431007374722e32002e4c706372656c5f6869333432002e4c706372656c5f6869333433002e4c616e6f6e2e31613066333665653566646430393230663564383432643039653237613465372e3439002e4c706372656c5f6869333439002e4c706372656c5f6869333538002e4c706372656c5f6869333539002e4c706372656c5f6869333639002e4c4a54493139315f30002e4c42423139315f333137002e4c42423139315f323530002e4c42423139315f323537002e4c42423139315f323631002e4c42423139315f323733002e4c42423139315f323739002e4c706372656c5f6869333436002e4c706372656c5f6869333438002e4c706372656c5f6869333631002e4c706372656c5f6869333632002e4c706372656c5f6869333633002e4c706372656c5f6869333735002e4c706372656c5f6869333733002e4c706372656c5f6869333630002e4c706372656c5f6869333634002e4c706372656c5f6869333635002e4c706372656c5f6869333636002e4c706372656c5f6869333531002e4c706372656c5f6869333532002e4c706372656c5f6869333435002e4c706372656c5f6869333437002e4c706372656c5f6869333637002e4c706372656c5f6869333638002e4c706372656c5f6869333530002e4c706372656c5f6869333536002e4c706372656c5f6869333537002e4c706372656c5f6869333533002e4c706372656c5f6869333534002e4c706372656c5f6869333535002e4c706372656c5f6869333731002e4c706372656c5f6869333732002e4c706372656c5f6869333730002e4c706372656c5f6869333736002e4c706372656c5f6869333734005f5a4e397374616b655f736d7431315f42554444595f484541503137686233373038373966306266356136656445005f5a4e397374616b655f736d7431375f46495845445f424c4f434b5f484541503137683263393037643763366462633565363545002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3134002e4c616e6f6e2e38303935383932396432623564383039666666643062303138613637613331642e3237002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3732002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3733002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3734002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3735002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3736002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3737002e4c616e6f6e2e38633938333365666432613364636138373061653139336163333463643164312e3738002e4c6c696e655f7461626c655f737461727430002e4c6c696e655f7461626c655f73746172743100626c616b6532622d7265662e63006c6f61643634002478007365637572655f7a65726f5f6d656d6f7279002478006d656d7365745f762e3000626c616b6532625f636f6d707265737300247800626c616b6532625f7570646174652e706172742e30002478002478002478002478002478002e4c3020002e4c3020002e4c3020002e4c3020002e4c3020002e4c3020002e4c3020002e4c3020002e4c3020002e4c34002e4c35002e4c3130002e4c3132002e4c3131002e4c3020002e4c3020002e4c3020002e4c3020002e4c3020002e4c3020002e4c3020002e4c3020002e4c3135002e4c3236002e4c3434002e4c3438002e4c3531002e4c3532006c69622e63002478002478002478002478002e4c32002e4c33002e4c3335002e4c3437002e4c3132002e4c3739002e4c3830002e4c3134002e4c3135002e4c3136002e4c3831002e4c3138002e4c3230002e4c3231002e4c3738002e4c3235002e4c3236002e4c3237002e4c3238002e4c3331002e4c3332002e4c3333002e4c3334002e4c3330002e4c3137002e4c3239002e4c3130002e4c313433002e4c313437002e4c313438002e4c313439002e4c323033002e4c313532002e4c323034002e4c313735002e4c313736002e4c313632002e4c323031002e4c313737002e4c313638002e4c313730002e4c313738002e4c313731002e4c313733002e4c313536002e4c313539002e4c313630002e4c313631002e4c313634002e4c323035002e4c313537002e4c313637002e4c313534005f5f636b625f7374645f6d61696e005f7374617274006d656d6d6f7665006d656d637079006d656d636d70006d656d73657400626c616b6532625f75706461746500626c616b6532625f66696e616c00626c616b6532625f696e69745f6b65795f776974685f706172616d00626c616b6532625f696e69745f706172616d000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001000000120000000000000060010100000000006001000000000000100d00000000000000000000000000001000000000000000000000000000000009000000010000001200000000000000700e010000000000700e000000000000400000000000000000000000000000000800000000000000080000000000000017000000010000000200000000000000b00e010000000000b00e000000000000c4170000000000000000000000000000080000000000000000000000000000002100000001000000060000000000000074360100000000007426000000000000be820100000000000000000000000000040000000000000000000000000000002700000001000000030000000000000038c902000000000038a9010000000000a8000000000000000000000000000000080000000000000000000000000000002e000000010000000300000000000000e0c9020000000000e0a9010000000000b8000000000000000000000000000000080000000000000000000000000000003400000001000000030000000000000098ca02000000000098aa010000000000080000000000000000000000000000000800000000000000000000000000000046000000080000000300000000000000a0ca020000000000a0aa01000000000000200800000000000000000000000000010000000000000000000000000000004b0000000100000000000000000000000000000000000000a0aa0100000000002802000000000000000000000000000001000000000000000000000000000000590000000100000000000000000000000000000000000000c8ac0100000000009c2600000000000000000000000000000100000000000000000000000000000065000000010000000000000000000000000000000000000064d3010000000000300200000000000000000000000000000100000000000000000000000000000074000000010000000000000000000000000000000000000094d5010000000000801300000000000000000000000000000100000000000000000000000000000082000000010000003000000000000000000000000000000014e901000000000012500000000000000000000000000000010000000000000001000000000000008d000000010000000000000000000000000000000000000026390200000000005d1c0000000000000000000000000000010000000000000000000000000000009d000000010000000000000000000000000000000000000083550200000000002400000000000000000000000000000001000000000000000000000000000000ad0000000300007000000000000000000000000000000000a7550200000000002b00000000000000000000000000000001000000000000000000000000000000bf0000000100000000000000000000000000000000000000d255020000000000041f000000000000000000000000000001000000000000000000000000000000cb0000000100000030000000000000000000000000000000d6740200000000002300000000000000000000000000000001000000000000000100000000000000d400000002000000000000000000000000000000000000000075020000000000c82d010000000000150000008d0c000008000000000000001800000000000000dc0000000300000000000000000000000000000000000000c8a2030000000000ee00000000000000000000000000000001000000000000000000000000000000e60000000300000000000000000000000000000000000000b6a3030000000000086c000000000000000000000000000001000000000000000000000000000000",
      "0x"
    ],
    "witnesses": [
      "0x55000000100000005500000055000000410000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
      "0x"
    ]
  },
  "cell_tx_signatures": {
    "0x61a0d1fa2b4a4536a778659d5d87b88e82188b17": [
      "0x861cb49aeea4929ad8af72e33591ec1db7330103907b084a9d6d3e507698d79819de6584720f26e961022e25a0efc9ef6a26ff9fa58c954dfd6989f9c5db4be400"
    ]
  },
  "cell_changes": [
    {
      "name": "stake",
      "kind": "NewAdded",
      "old_capacity": 0,
      "new_capacity": 16298200000000
    },
    {
      "name": "stake-smt",
      "kind": "NewAdded",
      "old_capacity": 0,
      "new_capacity": 26771000000000
    }
  ],
  "dep_group_tx": null,
  "dep_group_tx_signatures": {},
  "dep_group_changes": []
}